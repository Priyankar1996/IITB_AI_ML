-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_34_start: Boolean;
  signal convTranspose_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_540_inst_req_1 : boolean;
  signal type_cast_598_inst_ack_0 : boolean;
  signal type_cast_733_inst_req_0 : boolean;
  signal WPIPE_Block0_start_985_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_ack_1 : boolean;
  signal type_cast_598_inst_req_0 : boolean;
  signal addr_of_695_final_reg_req_1 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1085_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1064_inst_ack_0 : boolean;
  signal type_cast_733_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1003_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_ack_1 : boolean;
  signal type_cast_544_inst_ack_1 : boolean;
  signal type_cast_544_inst_req_1 : boolean;
  signal type_cast_598_inst_ack_1 : boolean;
  signal type_cast_544_inst_ack_0 : boolean;
  signal type_cast_544_inst_req_0 : boolean;
  signal type_cast_598_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1044_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_ack_1 : boolean;
  signal addr_of_695_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_req_1 : boolean;
  signal type_cast_45_inst_req_0 : boolean;
  signal type_cast_45_inst_ack_0 : boolean;
  signal type_cast_45_inst_req_1 : boolean;
  signal type_cast_45_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1044_inst_ack_0 : boolean;
  signal type_cast_1411_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_54_inst_ack_1 : boolean;
  signal type_cast_715_inst_ack_0 : boolean;
  signal if_stmt_638_branch_req_0 : boolean;
  signal type_cast_58_inst_req_0 : boolean;
  signal type_cast_58_inst_ack_0 : boolean;
  signal type_cast_58_inst_req_1 : boolean;
  signal type_cast_58_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1017_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_1 : boolean;
  signal ptr_deref_624_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1070_inst_req_1 : boolean;
  signal addr_of_695_final_reg_req_0 : boolean;
  signal type_cast_715_inst_req_0 : boolean;
  signal type_cast_70_inst_req_0 : boolean;
  signal type_cast_70_inst_ack_0 : boolean;
  signal array_obj_ref_694_index_offset_ack_1 : boolean;
  signal type_cast_70_inst_req_1 : boolean;
  signal ptr_deref_624_store_0_req_1 : boolean;
  signal type_cast_70_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_594_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1064_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_79_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1070_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_req_1 : boolean;
  signal array_obj_ref_694_index_offset_req_1 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_req_0 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_req_1 : boolean;
  signal type_cast_665_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1017_inst_req_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal type_cast_1401_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_ack_0 : boolean;
  signal type_cast_665_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_104_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_ack_0 : boolean;
  signal type_cast_616_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1064_inst_ack_1 : boolean;
  signal type_cast_108_inst_req_0 : boolean;
  signal type_cast_108_inst_ack_0 : boolean;
  signal array_obj_ref_694_index_offset_ack_0 : boolean;
  signal type_cast_108_inst_req_1 : boolean;
  signal ptr_deref_624_store_0_ack_0 : boolean;
  signal type_cast_108_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1003_inst_req_0 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_0 : boolean;
  signal type_cast_665_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 : boolean;
  signal type_cast_580_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_1 : boolean;
  signal ptr_deref_624_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_req_0 : boolean;
  signal type_cast_616_inst_req_1 : boolean;
  signal type_cast_120_inst_req_0 : boolean;
  signal type_cast_120_inst_ack_0 : boolean;
  signal array_obj_ref_694_index_offset_req_0 : boolean;
  signal type_cast_120_inst_req_1 : boolean;
  signal type_cast_120_inst_ack_1 : boolean;
  signal type_cast_715_inst_ack_1 : boolean;
  signal type_cast_733_inst_ack_1 : boolean;
  signal type_cast_580_inst_req_1 : boolean;
  signal type_cast_665_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_129_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1017_inst_ack_1 : boolean;
  signal type_cast_133_inst_req_0 : boolean;
  signal type_cast_133_inst_ack_0 : boolean;
  signal type_cast_133_inst_req_1 : boolean;
  signal type_cast_133_inst_ack_1 : boolean;
  signal type_cast_715_inst_req_1 : boolean;
  signal type_cast_733_inst_req_1 : boolean;
  signal type_cast_1401_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 : boolean;
  signal type_cast_580_inst_ack_0 : boolean;
  signal type_cast_346_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1020_inst_ack_0 : boolean;
  signal type_cast_346_inst_ack_0 : boolean;
  signal type_cast_346_inst_req_1 : boolean;
  signal type_cast_346_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_355_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_0 : boolean;
  signal type_cast_145_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_1 : boolean;
  signal type_cast_145_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_0 : boolean;
  signal type_cast_580_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_698_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_154_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_ack_0 : boolean;
  signal type_cast_616_inst_ack_0 : boolean;
  signal type_cast_158_inst_req_0 : boolean;
  signal type_cast_158_inst_ack_0 : boolean;
  signal type_cast_158_inst_req_1 : boolean;
  signal type_cast_158_inst_ack_1 : boolean;
  signal addr_of_695_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1044_inst_req_0 : boolean;
  signal type_cast_170_inst_req_0 : boolean;
  signal type_cast_170_inst_ack_0 : boolean;
  signal type_cast_170_inst_req_1 : boolean;
  signal type_cast_170_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1076_inst_ack_0 : boolean;
  signal type_cast_616_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_179_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_ack_0 : boolean;
  signal type_cast_183_inst_req_0 : boolean;
  signal type_cast_183_inst_ack_0 : boolean;
  signal type_cast_183_inst_req_1 : boolean;
  signal type_cast_183_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_576_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_979_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_576_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_ack_1 : boolean;
  signal type_cast_702_inst_ack_1 : boolean;
  signal type_cast_702_inst_req_1 : boolean;
  signal WPIPE_Block0_start_988_inst_req_0 : boolean;
  signal type_cast_195_inst_req_0 : boolean;
  signal type_cast_195_inst_ack_0 : boolean;
  signal type_cast_195_inst_req_1 : boolean;
  signal type_cast_195_inst_ack_1 : boolean;
  signal if_stmt_638_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1044_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_204_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_204_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_576_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_204_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_204_inst_ack_1 : boolean;
  signal type_cast_208_inst_req_0 : boolean;
  signal type_cast_208_inst_ack_0 : boolean;
  signal type_cast_208_inst_req_1 : boolean;
  signal type_cast_208_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_576_inst_req_0 : boolean;
  signal type_cast_217_inst_req_0 : boolean;
  signal type_cast_217_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_req_0 : boolean;
  signal type_cast_217_inst_req_1 : boolean;
  signal type_cast_217_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal type_cast_221_inst_req_0 : boolean;
  signal type_cast_221_inst_ack_0 : boolean;
  signal type_cast_221_inst_req_1 : boolean;
  signal type_cast_221_inst_ack_1 : boolean;
  signal type_cast_1055_inst_ack_0 : boolean;
  signal type_cast_225_inst_req_0 : boolean;
  signal type_cast_225_inst_ack_0 : boolean;
  signal type_cast_225_inst_req_1 : boolean;
  signal type_cast_225_inst_ack_1 : boolean;
  signal type_cast_562_inst_ack_1 : boolean;
  signal type_cast_562_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_req_1 : boolean;
  signal type_cast_262_inst_req_0 : boolean;
  signal type_cast_262_inst_ack_0 : boolean;
  signal type_cast_262_inst_req_1 : boolean;
  signal type_cast_262_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_0 : boolean;
  signal type_cast_266_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_1 : boolean;
  signal type_cast_266_inst_ack_1 : boolean;
  signal type_cast_562_inst_ack_0 : boolean;
  signal type_cast_562_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_612_inst_req_0 : boolean;
  signal type_cast_270_inst_req_0 : boolean;
  signal type_cast_270_inst_ack_0 : boolean;
  signal type_cast_270_inst_req_1 : boolean;
  signal type_cast_270_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1017_inst_ack_0 : boolean;
  signal type_cast_274_inst_req_0 : boolean;
  signal type_cast_274_inst_ack_0 : boolean;
  signal type_cast_274_inst_req_1 : boolean;
  signal type_cast_274_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_292_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_292_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_292_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_292_inst_ack_1 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal type_cast_296_inst_req_0 : boolean;
  signal type_cast_296_inst_ack_0 : boolean;
  signal type_cast_296_inst_req_1 : boolean;
  signal type_cast_296_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_558_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_558_inst_req_1 : boolean;
  signal WPIPE_Block0_start_979_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_req_0 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_305_inst_ack_1 : boolean;
  signal type_cast_702_inst_ack_0 : boolean;
  signal type_cast_702_inst_req_0 : boolean;
  signal type_cast_309_inst_req_0 : boolean;
  signal type_cast_309_inst_ack_0 : boolean;
  signal type_cast_309_inst_req_1 : boolean;
  signal type_cast_309_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_558_inst_ack_0 : boolean;
  signal if_stmt_638_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_558_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_317_inst_ack_1 : boolean;
  signal type_cast_321_inst_req_0 : boolean;
  signal WPIPE_Block0_start_988_inst_req_1 : boolean;
  signal type_cast_321_inst_ack_0 : boolean;
  signal type_cast_321_inst_req_1 : boolean;
  signal type_cast_321_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_330_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_330_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_330_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_330_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_req_0 : boolean;
  signal type_cast_334_inst_req_0 : boolean;
  signal type_cast_334_inst_ack_0 : boolean;
  signal type_cast_334_inst_req_1 : boolean;
  signal type_cast_334_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_342_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_342_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_342_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_342_inst_ack_1 : boolean;
  signal type_cast_359_inst_req_0 : boolean;
  signal type_cast_359_inst_ack_0 : boolean;
  signal type_cast_359_inst_req_1 : boolean;
  signal type_cast_359_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1003_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_367_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1003_inst_ack_1 : boolean;
  signal type_cast_1401_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1020_inst_req_1 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_380_inst_req_0 : boolean;
  signal WPIPE_Block0_start_997_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_380_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_380_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_380_inst_ack_1 : boolean;
  signal type_cast_1289_inst_ack_1 : boolean;
  signal type_cast_1401_inst_req_1 : boolean;
  signal type_cast_384_inst_req_0 : boolean;
  signal type_cast_384_inst_ack_0 : boolean;
  signal type_cast_384_inst_req_1 : boolean;
  signal type_cast_384_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_392_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_392_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_392_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_392_inst_ack_1 : boolean;
  signal type_cast_396_inst_req_0 : boolean;
  signal type_cast_396_inst_ack_0 : boolean;
  signal type_cast_396_inst_req_1 : boolean;
  signal type_cast_396_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_405_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_405_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_405_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_405_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1023_inst_req_1 : boolean;
  signal type_cast_409_inst_req_0 : boolean;
  signal type_cast_409_inst_ack_0 : boolean;
  signal type_cast_409_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_ack_1 : boolean;
  signal type_cast_409_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_req_0 : boolean;
  signal WPIPE_Block0_start_982_inst_req_0 : boolean;
  signal if_stmt_422_branch_req_0 : boolean;
  signal if_stmt_422_branch_ack_1 : boolean;
  signal if_stmt_422_branch_ack_0 : boolean;
  signal if_stmt_437_branch_req_0 : boolean;
  signal if_stmt_437_branch_ack_1 : boolean;
  signal if_stmt_437_branch_ack_0 : boolean;
  signal type_cast_458_inst_req_0 : boolean;
  signal type_cast_458_inst_ack_0 : boolean;
  signal type_cast_458_inst_req_1 : boolean;
  signal type_cast_458_inst_ack_1 : boolean;
  signal array_obj_ref_487_index_offset_req_0 : boolean;
  signal array_obj_ref_487_index_offset_ack_0 : boolean;
  signal array_obj_ref_487_index_offset_req_1 : boolean;
  signal array_obj_ref_487_index_offset_ack_1 : boolean;
  signal addr_of_488_final_reg_req_0 : boolean;
  signal addr_of_488_final_reg_ack_0 : boolean;
  signal addr_of_488_final_reg_req_1 : boolean;
  signal addr_of_488_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_491_inst_ack_1 : boolean;
  signal type_cast_495_inst_req_0 : boolean;
  signal type_cast_495_inst_ack_0 : boolean;
  signal type_cast_495_inst_req_1 : boolean;
  signal type_cast_495_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_ack_1 : boolean;
  signal type_cast_508_inst_req_0 : boolean;
  signal type_cast_508_inst_ack_0 : boolean;
  signal type_cast_508_inst_req_1 : boolean;
  signal type_cast_508_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_ack_1 : boolean;
  signal type_cast_526_inst_req_0 : boolean;
  signal type_cast_526_inst_ack_0 : boolean;
  signal type_cast_526_inst_req_1 : boolean;
  signal type_cast_526_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1064_inst_req_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_req_1 : boolean;
  signal type_cast_1411_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_765_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1041_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_765_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_765_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1041_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_765_inst_ack_1 : boolean;
  signal type_cast_769_inst_req_0 : boolean;
  signal type_cast_769_inst_ack_0 : boolean;
  signal type_cast_769_inst_req_1 : boolean;
  signal type_cast_769_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_783_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1041_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_783_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_783_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1041_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_783_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1014_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1014_inst_req_1 : boolean;
  signal type_cast_787_inst_req_0 : boolean;
  signal type_cast_787_inst_ack_0 : boolean;
  signal type_cast_787_inst_req_1 : boolean;
  signal type_cast_787_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1082_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_801_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_801_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_991_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_801_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_801_inst_ack_1 : boolean;
  signal type_cast_805_inst_req_0 : boolean;
  signal type_cast_805_inst_ack_0 : boolean;
  signal type_cast_805_inst_req_1 : boolean;
  signal type_cast_805_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_819_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_819_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_991_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_819_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_819_inst_ack_1 : boolean;
  signal if_stmt_1316_branch_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1014_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1014_inst_req_0 : boolean;
  signal type_cast_823_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_req_1 : boolean;
  signal type_cast_823_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1073_inst_ack_1 : boolean;
  signal type_cast_823_inst_req_1 : boolean;
  signal type_cast_823_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1038_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_req_0 : boolean;
  signal ptr_deref_831_store_0_req_0 : boolean;
  signal ptr_deref_831_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_req_1 : boolean;
  signal ptr_deref_831_store_0_req_1 : boolean;
  signal ptr_deref_831_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1073_inst_req_1 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_0 : boolean;
  signal if_stmt_845_branch_req_0 : boolean;
  signal WPIPE_Block0_start_985_inst_req_0 : boolean;
  signal if_stmt_845_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1029_inst_ack_0 : boolean;
  signal if_stmt_845_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1070_inst_ack_0 : boolean;
  signal type_cast_856_inst_req_0 : boolean;
  signal type_cast_856_inst_ack_0 : boolean;
  signal type_cast_856_inst_req_1 : boolean;
  signal type_cast_856_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1079_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1076_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1073_inst_ack_0 : boolean;
  signal type_cast_860_inst_req_0 : boolean;
  signal type_cast_860_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1073_inst_req_0 : boolean;
  signal type_cast_860_inst_req_1 : boolean;
  signal type_cast_860_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1079_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_ack_1 : boolean;
  signal type_cast_1062_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_req_0 : boolean;
  signal type_cast_1343_inst_req_0 : boolean;
  signal type_cast_864_inst_req_0 : boolean;
  signal type_cast_864_inst_ack_0 : boolean;
  signal type_cast_864_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_ack_1 : boolean;
  signal type_cast_864_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_req_0 : boolean;
  signal if_stmt_882_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1011_inst_req_0 : boolean;
  signal if_stmt_882_branch_ack_1 : boolean;
  signal if_stmt_882_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_ack_1 : boolean;
  signal type_cast_1062_inst_req_1 : boolean;
  signal type_cast_909_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1035_inst_req_1 : boolean;
  signal type_cast_909_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_req_1 : boolean;
  signal type_cast_909_inst_req_1 : boolean;
  signal type_cast_909_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1070_inst_req_0 : boolean;
  signal type_cast_1062_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_1 : boolean;
  signal if_stmt_1316_branch_ack_0 : boolean;
  signal array_obj_ref_938_index_offset_req_0 : boolean;
  signal array_obj_ref_938_index_offset_ack_0 : boolean;
  signal array_obj_ref_938_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_ack_0 : boolean;
  signal array_obj_ref_938_index_offset_ack_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_req_0 : boolean;
  signal addr_of_939_final_reg_req_0 : boolean;
  signal addr_of_939_final_reg_ack_0 : boolean;
  signal addr_of_939_final_reg_req_1 : boolean;
  signal addr_of_939_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_req_0 : boolean;
  signal type_cast_1062_inst_req_0 : boolean;
  signal type_cast_1343_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1026_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1000_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_req_1 : boolean;
  signal ptr_deref_942_store_0_req_0 : boolean;
  signal ptr_deref_942_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_req_0 : boolean;
  signal WPIPE_Block0_start_982_inst_req_1 : boolean;
  signal ptr_deref_942_store_0_req_1 : boolean;
  signal ptr_deref_942_store_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1007_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1007_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_req_1 : boolean;
  signal if_stmt_957_branch_req_0 : boolean;
  signal if_stmt_957_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_0 : boolean;
  signal if_stmt_957_branch_ack_0 : boolean;
  signal call_stmt_968_call_req_0 : boolean;
  signal WPIPE_Block1_start_1032_inst_req_1 : boolean;
  signal call_stmt_968_call_ack_0 : boolean;
  signal type_cast_1343_inst_ack_0 : boolean;
  signal call_stmt_968_call_req_1 : boolean;
  signal call_stmt_968_call_ack_1 : boolean;
  signal type_cast_973_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1032_inst_ack_0 : boolean;
  signal type_cast_973_inst_ack_0 : boolean;
  signal type_cast_973_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_req_0 : boolean;
  signal type_cast_973_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_991_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_991_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1 : boolean;
  signal type_cast_1289_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1 : boolean;
  signal type_cast_1343_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_976_inst_req_0 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_0 : boolean;
  signal type_cast_1381_inst_req_0 : boolean;
  signal WPIPE_Block0_start_976_inst_req_1 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1094_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1094_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1097_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1097_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1097_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1097_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_ack_1 : boolean;
  signal ptr_deref_1377_load_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1100_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1300_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1100_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_req_1 : boolean;
  signal ptr_deref_1377_load_0_req_1 : boolean;
  signal if_stmt_1316_branch_req_0 : boolean;
  signal type_cast_1111_inst_req_0 : boolean;
  signal type_cast_1111_inst_ack_0 : boolean;
  signal type_cast_1111_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_ack_0 : boolean;
  signal type_cast_1411_inst_ack_0 : boolean;
  signal type_cast_1118_inst_req_0 : boolean;
  signal type_cast_1118_inst_ack_0 : boolean;
  signal type_cast_1411_inst_req_0 : boolean;
  signal type_cast_1118_inst_req_1 : boolean;
  signal type_cast_1118_inst_ack_1 : boolean;
  signal ptr_deref_1377_load_0_ack_0 : boolean;
  signal type_cast_1391_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1120_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1120_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1120_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1120_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1453_inst_req_0 : boolean;
  signal ptr_deref_1377_load_0_req_0 : boolean;
  signal type_cast_1391_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1123_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_req_1 : boolean;
  signal addr_of_1373_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1123_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1456_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1126_inst_req_0 : boolean;
  signal addr_of_1373_final_reg_req_1 : boolean;
  signal WPIPE_Block2_start_1126_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1126_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1126_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1312_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1129_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1129_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1129_inst_req_1 : boolean;
  signal addr_of_1373_final_reg_ack_0 : boolean;
  signal WPIPE_Block2_start_1129_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1459_inst_req_0 : boolean;
  signal type_cast_1451_inst_ack_1 : boolean;
  signal type_cast_1451_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1312_inst_req_1 : boolean;
  signal type_cast_1391_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_req_0 : boolean;
  signal addr_of_1373_final_reg_req_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1132_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1132_inst_ack_1 : boolean;
  signal type_cast_1391_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1135_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1135_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_ack_1 : boolean;
  signal type_cast_1451_inst_ack_0 : boolean;
  signal type_cast_1451_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1312_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1138_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1312_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1297_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_req_1 : boolean;
  signal array_obj_ref_1372_index_offset_ack_1 : boolean;
  signal WPIPE_Block3_start_1141_inst_ack_1 : boolean;
  signal type_cast_1441_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1144_inst_req_0 : boolean;
  signal array_obj_ref_1372_index_offset_req_1 : boolean;
  signal WPIPE_Block3_start_1144_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1144_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1144_inst_ack_1 : boolean;
  signal type_cast_1441_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1147_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1147_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_ack_1 : boolean;
  signal type_cast_1441_inst_ack_0 : boolean;
  signal type_cast_1441_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1150_inst_req_0 : boolean;
  signal array_obj_ref_1372_index_offset_ack_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_req_1 : boolean;
  signal array_obj_ref_1372_index_offset_req_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1153_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1153_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1153_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1153_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_1 : boolean;
  signal type_cast_1431_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_ack_0 : boolean;
  signal type_cast_1381_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1156_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1156_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1156_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1156_inst_ack_1 : boolean;
  signal type_cast_1431_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1309_inst_req_0 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_0 : boolean;
  signal type_cast_1381_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_1 : boolean;
  signal type_cast_1431_inst_ack_0 : boolean;
  signal type_cast_1431_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_req_1 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal type_cast_1174_inst_req_1 : boolean;
  signal type_cast_1174_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1176_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1176_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1306_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1179_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 : boolean;
  signal type_cast_1421_inst_ack_1 : boolean;
  signal type_cast_1421_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1182_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1182_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1182_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1182_inst_ack_1 : boolean;
  signal type_cast_1421_inst_ack_0 : boolean;
  signal type_cast_1381_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1185_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1185_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1185_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1185_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 : boolean;
  signal type_cast_1421_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1190_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1190_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1190_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1190_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1193_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1193_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1193_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1193_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1196_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1196_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1196_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1196_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1199_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1199_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1199_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1199_inst_ack_1 : boolean;
  signal call_stmt_1203_call_req_0 : boolean;
  signal call_stmt_1203_call_ack_0 : boolean;
  signal call_stmt_1203_call_req_1 : boolean;
  signal call_stmt_1203_call_ack_1 : boolean;
  signal type_cast_1207_inst_req_0 : boolean;
  signal type_cast_1207_inst_ack_0 : boolean;
  signal type_cast_1207_inst_req_1 : boolean;
  signal type_cast_1207_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1214_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1214_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1214_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1214_inst_ack_1 : boolean;
  signal type_cast_1219_inst_req_0 : boolean;
  signal type_cast_1219_inst_ack_0 : boolean;
  signal type_cast_1219_inst_req_1 : boolean;
  signal type_cast_1219_inst_ack_1 : boolean;
  signal type_cast_1229_inst_req_0 : boolean;
  signal type_cast_1229_inst_ack_0 : boolean;
  signal type_cast_1229_inst_req_1 : boolean;
  signal type_cast_1229_inst_ack_1 : boolean;
  signal type_cast_1239_inst_req_0 : boolean;
  signal type_cast_1239_inst_ack_0 : boolean;
  signal type_cast_1239_inst_req_1 : boolean;
  signal type_cast_1239_inst_ack_1 : boolean;
  signal type_cast_1249_inst_req_0 : boolean;
  signal type_cast_1249_inst_ack_0 : boolean;
  signal type_cast_1249_inst_req_1 : boolean;
  signal type_cast_1249_inst_ack_1 : boolean;
  signal type_cast_1259_inst_req_0 : boolean;
  signal type_cast_1259_inst_ack_0 : boolean;
  signal type_cast_1259_inst_req_1 : boolean;
  signal type_cast_1259_inst_ack_1 : boolean;
  signal type_cast_1269_inst_req_0 : boolean;
  signal type_cast_1269_inst_ack_0 : boolean;
  signal type_cast_1269_inst_req_1 : boolean;
  signal type_cast_1269_inst_ack_1 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal type_cast_1289_inst_req_0 : boolean;
  signal type_cast_1289_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1462_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1465_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1468_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1471_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1471_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1471_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1471_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1474_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1474_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1474_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1474_inst_ack_1 : boolean;
  signal if_stmt_1488_branch_req_0 : boolean;
  signal if_stmt_1488_branch_ack_1 : boolean;
  signal if_stmt_1488_branch_ack_0 : boolean;
  signal phi_stmt_475_req_0 : boolean;
  signal type_cast_481_inst_req_0 : boolean;
  signal type_cast_481_inst_ack_0 : boolean;
  signal type_cast_481_inst_req_1 : boolean;
  signal type_cast_481_inst_ack_1 : boolean;
  signal phi_stmt_475_req_1 : boolean;
  signal phi_stmt_475_ack_0 : boolean;
  signal phi_stmt_682_req_1 : boolean;
  signal type_cast_685_inst_req_0 : boolean;
  signal type_cast_685_inst_ack_0 : boolean;
  signal type_cast_685_inst_req_1 : boolean;
  signal type_cast_685_inst_ack_1 : boolean;
  signal phi_stmt_682_req_0 : boolean;
  signal phi_stmt_682_ack_0 : boolean;
  signal phi_stmt_926_req_1 : boolean;
  signal type_cast_929_inst_req_0 : boolean;
  signal type_cast_929_inst_ack_0 : boolean;
  signal type_cast_929_inst_req_1 : boolean;
  signal type_cast_929_inst_ack_1 : boolean;
  signal phi_stmt_926_req_0 : boolean;
  signal phi_stmt_926_ack_0 : boolean;
  signal phi_stmt_1360_req_0 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal phi_stmt_1360_req_1 : boolean;
  signal phi_stmt_1360_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_34: Block -- control-path 
    signal convTranspose_CP_34_elements: BooleanArray(500 downto 0);
    -- 
  begin -- 
    convTranspose_CP_34_elements(0) <= convTranspose_CP_34_start;
    convTranspose_CP_34_symbol <= convTranspose_CP_34_elements(500);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_39/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/branch_block_stmt_39__entry__
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421__entry__
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_update_start_
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Update/cr
      -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => RPIPE_ConvTranspose_input_pipe_41_inst_req_0); -- 
    cr_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_45_inst_req_1); -- 
    cr_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_58_inst_req_1); -- 
    cr_207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_70_inst_req_1); -- 
    cr_235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_83_inst_req_1); -- 
    cr_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_95_inst_req_1); -- 
    cr_291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_108_inst_req_1); -- 
    cr_319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_120_inst_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_133_inst_req_1); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_346_inst_req_1); -- 
    cr_375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_145_inst_req_1); -- 
    cr_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_158_inst_req_1); -- 
    cr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_170_inst_req_1); -- 
    cr_459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_183_inst_req_1); -- 
    cr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_195_inst_req_1); -- 
    cr_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_208_inst_req_1); -- 
    cr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_217_inst_req_1); -- 
    cr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_221_inst_req_1); -- 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_225_inst_req_1); -- 
    cr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_262_inst_req_1); -- 
    cr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_266_inst_req_1); -- 
    cr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_270_inst_req_1); -- 
    cr_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_274_inst_req_1); -- 
    cr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_296_inst_req_1); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_309_inst_req_1); -- 
    cr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_321_inst_req_1); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_334_inst_req_1); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_359_inst_req_1); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_371_inst_req_1); -- 
    cr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_384_inst_req_1); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_396_inst_req_1); -- 
    cr_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_409_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_update_start_
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Update/cr
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_41_inst_ack_0, ack => convTranspose_CP_34_elements(1)); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(1), ack => RPIPE_ConvTranspose_input_pipe_41_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_41_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_sample_start_
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_41_inst_ack_1, ack => convTranspose_CP_34_elements(2)); -- 
    rr_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => type_cast_45_inst_req_0); -- 
    rr_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => RPIPE_ConvTranspose_input_pipe_54_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Sample/ra
      -- 
    ra_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_0, ack => convTranspose_CP_34_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_45_Update/ca
      -- 
    ca_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_1, ack => convTranspose_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_update_start_
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Update/cr
      -- 
    ra_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_54_inst_ack_0, ack => convTranspose_CP_34_elements(5)); -- 
    cr_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(5), ack => RPIPE_ConvTranspose_input_pipe_54_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_54_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Sample/rr
      -- 
    ca_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_54_inst_ack_1, ack => convTranspose_CP_34_elements(6)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => type_cast_58_inst_req_0); -- 
    rr_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Sample/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_0, ack => convTranspose_CP_34_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_58_Update/ca
      -- 
    ca_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_58_inst_ack_1, ack => convTranspose_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_update_start_
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Update/cr
      -- 
    ra_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_0, ack => convTranspose_CP_34_elements(9)); -- 
    cr_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(9), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_66_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Sample/rr
      -- 
    ca_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_1, ack => convTranspose_CP_34_elements(10)); -- 
    rr_202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => type_cast_70_inst_req_0); -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => RPIPE_ConvTranspose_input_pipe_79_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Sample/ra
      -- 
    ra_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_0, ack => convTranspose_CP_34_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_70_Update/ca
      -- 
    ca_208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_1, ack => convTranspose_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_update_start_
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Update/cr
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_79_inst_ack_0, ack => convTranspose_CP_34_elements(13)); -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(13), ack => RPIPE_ConvTranspose_input_pipe_79_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_79_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Sample/rr
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_79_inst_ack_1, ack => convTranspose_CP_34_elements(14)); -- 
    rr_230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => type_cast_83_inst_req_0); -- 
    rr_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Sample/ra
      -- 
    ra_231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => convTranspose_CP_34_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_83_Update/ca
      -- 
    ca_236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => convTranspose_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_update_start_
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Update/cr
      -- 
    ra_245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_0, ack => convTranspose_CP_34_elements(17)); -- 
    cr_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(17), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_91_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Sample/rr
      -- 
    ca_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_1, ack => convTranspose_CP_34_elements(18)); -- 
    rr_258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => type_cast_95_inst_req_0); -- 
    rr_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => RPIPE_ConvTranspose_input_pipe_104_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Sample/ra
      -- 
    ra_259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => convTranspose_CP_34_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_95_Update/ca
      -- 
    ca_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => convTranspose_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_update_start_
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Update/cr
      -- 
    ra_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_104_inst_ack_0, ack => convTranspose_CP_34_elements(21)); -- 
    cr_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(21), ack => RPIPE_ConvTranspose_input_pipe_104_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_104_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Sample/rr
      -- 
    ca_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_104_inst_ack_1, ack => convTranspose_CP_34_elements(22)); -- 
    rr_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => type_cast_108_inst_req_0); -- 
    rr_300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Sample/ra
      -- 
    ra_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_0, ack => convTranspose_CP_34_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_108_Update/ca
      -- 
    ca_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_1, ack => convTranspose_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_update_start_
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Update/cr
      -- 
    ra_301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_0, ack => convTranspose_CP_34_elements(25)); -- 
    cr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(25), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_116_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Sample/rr
      -- 
    ca_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_1, ack => convTranspose_CP_34_elements(26)); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => type_cast_120_inst_req_0); -- 
    rr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => RPIPE_ConvTranspose_input_pipe_129_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Sample/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_0, ack => convTranspose_CP_34_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_120_Update/ca
      -- 
    ca_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_1, ack => convTranspose_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_update_start_
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Update/cr
      -- 
    ra_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_129_inst_ack_0, ack => convTranspose_CP_34_elements(29)); -- 
    cr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(29), ack => RPIPE_ConvTranspose_input_pipe_129_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_129_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Sample/rr
      -- 
    ca_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_129_inst_ack_1, ack => convTranspose_CP_34_elements(30)); -- 
    rr_342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => type_cast_133_inst_req_0); -- 
    rr_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Sample/ra
      -- 
    ra_343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_133_inst_ack_0, ack => convTranspose_CP_34_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_133_Update/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_133_inst_ack_1, ack => convTranspose_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_update_start_
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Sample/ra
      -- 
    ra_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_0, ack => convTranspose_CP_34_elements(33)); -- 
    cr_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(33), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_141_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Sample/rr
      -- 
    ca_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_1, ack => convTranspose_CP_34_elements(34)); -- 
    rr_370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => type_cast_145_inst_req_0); -- 
    rr_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => RPIPE_ConvTranspose_input_pipe_154_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Sample/ra
      -- 
    ra_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_0, ack => convTranspose_CP_34_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_145_Update/ca
      -- 
    ca_376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_1, ack => convTranspose_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_update_start_
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Update/cr
      -- 
    ra_385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_154_inst_ack_0, ack => convTranspose_CP_34_elements(37)); -- 
    cr_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(37), ack => RPIPE_ConvTranspose_input_pipe_154_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_154_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Sample/rr
      -- 
    ca_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_154_inst_ack_1, ack => convTranspose_CP_34_elements(38)); -- 
    rr_398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => type_cast_158_inst_req_0); -- 
    rr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Sample/ra
      -- 
    ra_399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_158_inst_ack_0, ack => convTranspose_CP_34_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_158_Update/ca
      -- 
    ca_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_158_inst_ack_1, ack => convTranspose_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_update_start_
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Update/cr
      -- 
    ra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_0, ack => convTranspose_CP_34_elements(41)); -- 
    cr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(41), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_166_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Sample/rr
      -- 
    ca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_1, ack => convTranspose_CP_34_elements(42)); -- 
    rr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => type_cast_170_inst_req_0); -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => RPIPE_ConvTranspose_input_pipe_179_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Sample/ra
      -- 
    ra_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_0, ack => convTranspose_CP_34_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_170_Update/ca
      -- 
    ca_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_1, ack => convTranspose_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_update_start_
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Update/cr
      -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_179_inst_ack_0, ack => convTranspose_CP_34_elements(45)); -- 
    cr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(45), ack => RPIPE_ConvTranspose_input_pipe_179_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_179_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Sample/rr
      -- 
    ca_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_179_inst_ack_1, ack => convTranspose_CP_34_elements(46)); -- 
    rr_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => type_cast_183_inst_req_0); -- 
    rr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => RPIPE_ConvTranspose_input_pipe_191_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Sample/ra
      -- 
    ra_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_183_inst_ack_0, ack => convTranspose_CP_34_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_183_Update/ca
      -- 
    ca_460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_183_inst_ack_1, ack => convTranspose_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_update_start_
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Update/cr
      -- 
    ra_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_191_inst_ack_0, ack => convTranspose_CP_34_elements(49)); -- 
    cr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(49), ack => RPIPE_ConvTranspose_input_pipe_191_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_191_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Sample/rr
      -- 
    ca_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_191_inst_ack_1, ack => convTranspose_CP_34_elements(50)); -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => type_cast_195_inst_req_0); -- 
    rr_496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => RPIPE_ConvTranspose_input_pipe_204_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Sample/ra
      -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_0, ack => convTranspose_CP_34_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_195_Update/ca
      -- 
    ca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_1, ack => convTranspose_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_update_start_
      -- CP-element group 53: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Update/cr
      -- 
    ra_497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_204_inst_ack_0, ack => convTranspose_CP_34_elements(53)); -- 
    cr_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(53), ack => RPIPE_ConvTranspose_input_pipe_204_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_204_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Sample/rr
      -- 
    ca_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_204_inst_ack_1, ack => convTranspose_CP_34_elements(54)); -- 
    rr_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => type_cast_208_inst_req_0); -- 
    rr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => RPIPE_ConvTranspose_input_pipe_292_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Sample/ra
      -- 
    ra_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_208_inst_ack_0, ack => convTranspose_CP_34_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_208_Update/ca
      -- 
    ca_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_208_inst_ack_1, ack => convTranspose_CP_34_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Sample/rr
      -- 
    rr_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(57), ack => type_cast_217_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(4) & convTranspose_CP_34_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Sample/ra
      -- 
    ra_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_217_inst_ack_0, ack => convTranspose_CP_34_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_217_Update/ca
      -- 
    ca_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_217_inst_ack_1, ack => convTranspose_CP_34_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Sample/rr
      -- 
    rr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(60), ack => type_cast_221_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(12) & convTranspose_CP_34_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Sample/ra
      -- 
    ra_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_221_inst_ack_0, ack => convTranspose_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_221_Update/ca
      -- 
    ca_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_221_inst_ack_1, ack => convTranspose_CP_34_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Sample/rr
      -- 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(63), ack => type_cast_225_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(20) & convTranspose_CP_34_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Sample/ra
      -- 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_225_inst_ack_0, ack => convTranspose_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_225_Update/ca
      -- 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_225_inst_ack_1, ack => convTranspose_CP_34_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Sample/rr
      -- 
    rr_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(66), ack => type_cast_262_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(28) & convTranspose_CP_34_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Sample/ra
      -- 
    ra_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_262_inst_ack_0, ack => convTranspose_CP_34_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_262_Update/ca
      -- 
    ca_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_262_inst_ack_1, ack => convTranspose_CP_34_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Sample/rr
      -- 
    rr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(69), ack => type_cast_266_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(40) & convTranspose_CP_34_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Sample/ra
      -- 
    ra_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_0, ack => convTranspose_CP_34_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_266_Update/ca
      -- 
    ca_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_1, ack => convTranspose_CP_34_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Sample/rr
      -- 
    rr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(72), ack => type_cast_270_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(44) & convTranspose_CP_34_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Sample/ra
      -- 
    ra_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_0, ack => convTranspose_CP_34_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_270_Update/ca
      -- 
    ca_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_1, ack => convTranspose_CP_34_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Sample/rr
      -- 
    rr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(75), ack => type_cast_274_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(52) & convTranspose_CP_34_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Sample/ra
      -- 
    ra_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_274_inst_ack_0, ack => convTranspose_CP_34_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_274_Update/ca
      -- 
    ca_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_274_inst_ack_1, ack => convTranspose_CP_34_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_update_start_
      -- CP-element group 78: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Update/cr
      -- 
    ra_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_292_inst_ack_0, ack => convTranspose_CP_34_elements(78)); -- 
    cr_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(78), ack => RPIPE_ConvTranspose_input_pipe_292_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_292_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Sample/rr
      -- 
    ca_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_292_inst_ack_1, ack => convTranspose_CP_34_elements(79)); -- 
    rr_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => type_cast_296_inst_req_0); -- 
    rr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => RPIPE_ConvTranspose_input_pipe_305_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Sample/ra
      -- 
    ra_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_296_inst_ack_0, ack => convTranspose_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_296_Update/ca
      -- 
    ca_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_296_inst_ack_1, ack => convTranspose_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_update_start_
      -- CP-element group 82: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Update/cr
      -- 
    ra_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_305_inst_ack_0, ack => convTranspose_CP_34_elements(82)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(82), ack => RPIPE_ConvTranspose_input_pipe_305_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_305_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Sample/rr
      -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_305_inst_ack_1, ack => convTranspose_CP_34_elements(83)); -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => type_cast_309_inst_req_0); -- 
    rr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => RPIPE_ConvTranspose_input_pipe_317_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Sample/ra
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_0, ack => convTranspose_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_309_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_1, ack => convTranspose_CP_34_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_update_start_
      -- CP-element group 86: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Update/cr
      -- 
    ra_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_317_inst_ack_0, ack => convTranspose_CP_34_elements(86)); -- 
    cr_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(86), ack => RPIPE_ConvTranspose_input_pipe_317_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_317_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Sample/rr
      -- 
    ca_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_317_inst_ack_1, ack => convTranspose_CP_34_elements(87)); -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => type_cast_321_inst_req_0); -- 
    rr_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => RPIPE_ConvTranspose_input_pipe_330_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Sample/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_321_inst_ack_0, ack => convTranspose_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_321_Update/ca
      -- 
    ca_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_321_inst_ack_1, ack => convTranspose_CP_34_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_update_start_
      -- CP-element group 90: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Update/cr
      -- 
    ra_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_330_inst_ack_0, ack => convTranspose_CP_34_elements(90)); -- 
    cr_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(90), ack => RPIPE_ConvTranspose_input_pipe_330_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_330_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Sample/rr
      -- 
    ca_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_330_inst_ack_1, ack => convTranspose_CP_34_elements(91)); -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => type_cast_334_inst_req_0); -- 
    rr_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => RPIPE_ConvTranspose_input_pipe_342_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Sample/ra
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_334_inst_ack_0, ack => convTranspose_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_334_Update/ca
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_334_inst_ack_1, ack => convTranspose_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_update_start_
      -- CP-element group 94: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Update/cr
      -- 
    ra_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_342_inst_ack_0, ack => convTranspose_CP_34_elements(94)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(94), ack => RPIPE_ConvTranspose_input_pipe_342_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_342_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Sample/$entry
      -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_342_inst_ack_1, ack => convTranspose_CP_34_elements(95)); -- 
    rr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => type_cast_346_inst_req_0); -- 
    rr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => RPIPE_ConvTranspose_input_pipe_355_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Sample/$exit
      -- 
    ra_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_346_inst_ack_0, ack => convTranspose_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_346_update_completed_
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_346_inst_ack_1, ack => convTranspose_CP_34_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_update_start_
      -- CP-element group 98: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Update/cr
      -- 
    ra_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_355_inst_ack_0, ack => convTranspose_CP_34_elements(98)); -- 
    cr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(98), ack => RPIPE_ConvTranspose_input_pipe_355_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_355_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Sample/rr
      -- 
    ca_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_355_inst_ack_1, ack => convTranspose_CP_34_elements(99)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => type_cast_359_inst_req_0); -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => RPIPE_ConvTranspose_input_pipe_367_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Sample/ra
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_0, ack => convTranspose_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_359_Update/ca
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_359_inst_ack_1, ack => convTranspose_CP_34_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_update_start_
      -- CP-element group 102: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Update/cr
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_367_inst_ack_0, ack => convTranspose_CP_34_elements(102)); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(102), ack => RPIPE_ConvTranspose_input_pipe_367_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_367_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Sample/rr
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_367_inst_ack_1, ack => convTranspose_CP_34_elements(103)); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => type_cast_371_inst_req_0); -- 
    rr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => RPIPE_ConvTranspose_input_pipe_380_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Sample/ra
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => convTranspose_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_371_Update/ca
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => convTranspose_CP_34_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_update_start_
      -- CP-element group 106: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Update/cr
      -- 
    ra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_380_inst_ack_0, ack => convTranspose_CP_34_elements(106)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(106), ack => RPIPE_ConvTranspose_input_pipe_380_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_380_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Sample/rr
      -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_380_inst_ack_1, ack => convTranspose_CP_34_elements(107)); -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => type_cast_384_inst_req_0); -- 
    rr_846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => RPIPE_ConvTranspose_input_pipe_392_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Sample/ra
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_384_inst_ack_0, ack => convTranspose_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_384_Update/ca
      -- 
    ca_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_384_inst_ack_1, ack => convTranspose_CP_34_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_update_start_
      -- CP-element group 110: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Update/cr
      -- 
    ra_847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_392_inst_ack_0, ack => convTranspose_CP_34_elements(110)); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(110), ack => RPIPE_ConvTranspose_input_pipe_392_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_392_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Sample/rr
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_392_inst_ack_1, ack => convTranspose_CP_34_elements(111)); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => type_cast_396_inst_req_0); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => RPIPE_ConvTranspose_input_pipe_405_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Sample/ra
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_396_inst_ack_0, ack => convTranspose_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_396_Update/ca
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_396_inst_ack_1, ack => convTranspose_CP_34_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_update_start_
      -- CP-element group 114: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Update/cr
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_405_inst_ack_0, ack => convTranspose_CP_34_elements(114)); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(114), ack => RPIPE_ConvTranspose_input_pipe_405_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/RPIPE_ConvTranspose_input_pipe_405_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Sample/rr
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_405_inst_ack_1, ack => convTranspose_CP_34_elements(115)); -- 
    rr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(115), ack => type_cast_409_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Sample/ra
      -- 
    ra_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_409_inst_ack_0, ack => convTranspose_CP_34_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/type_cast_409_Update/ca
      -- 
    ca_894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_409_inst_ack_1, ack => convTranspose_CP_34_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421__exit__
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422__entry__
      -- CP-element group 118: 	 branch_block_stmt_39/assign_stmt_42_to_assign_stmt_421/$exit
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_39/R_cmp514_423_place
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_39/if_stmt_422_else_link/$entry
      -- 
    branch_req_902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(118), ack => if_stmt_422_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(59) & convTranspose_CP_34_elements(62) & convTranspose_CP_34_elements(65) & convTranspose_CP_34_elements(68) & convTranspose_CP_34_elements(71) & convTranspose_CP_34_elements(74) & convTranspose_CP_34_elements(77) & convTranspose_CP_34_elements(81) & convTranspose_CP_34_elements(85) & convTranspose_CP_34_elements(89) & convTranspose_CP_34_elements(93) & convTranspose_CP_34_elements(97) & convTranspose_CP_34_elements(101) & convTranspose_CP_34_elements(105) & convTranspose_CP_34_elements(109) & convTranspose_CP_34_elements(113) & convTranspose_CP_34_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_39/merge_stmt_443__exit__
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472__entry__
      -- CP-element group 119: 	 branch_block_stmt_39/if_stmt_422_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_39/if_stmt_422_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_39/entry_bbx_xnph516
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/$entry
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_update_start_
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_39/entry_bbx_xnph516_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_39/entry_bbx_xnph516_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_39/merge_stmt_443_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_39/merge_stmt_443_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_39/merge_stmt_443_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_39/merge_stmt_443_PhiAck/dummy
      -- 
    if_choice_transition_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_422_branch_ack_1, ack => convTranspose_CP_34_elements(119)); -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_458_inst_req_0); -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_458_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	473 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_39/if_stmt_422_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_39/if_stmt_422_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_39/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_39/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_39/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_422_branch_ack_0, ack => convTranspose_CP_34_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	473 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_39/merge_stmt_644__exit__
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679__entry__
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_update_start_
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/$entry
      -- CP-element group 121: 	 branch_block_stmt_39/if_stmt_437_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_39/if_stmt_437_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_39/forx_xcond190x_xpreheader_bbx_xnph512
      -- CP-element group 121: 	 branch_block_stmt_39/forx_xcond190x_xpreheader_bbx_xnph512_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_39/forx_xcond190x_xpreheader_bbx_xnph512_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_39/merge_stmt_644_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_39/merge_stmt_644_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_39/merge_stmt_644_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_39/merge_stmt_644_PhiAck/dummy
      -- 
    if_choice_transition_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_437_branch_ack_1, ack => convTranspose_CP_34_elements(121)); -- 
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_665_inst_req_1); -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_665_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	473 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	486 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_39/if_stmt_437_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_39/if_stmt_437_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_39/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_39/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_39/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_437_branch_ack_0, ack => convTranspose_CP_34_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Sample/ra
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_0, ack => convTranspose_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	474 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472__exit__
      -- CP-element group 124: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/$exit
      -- CP-element group 124: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_39/assign_stmt_449_to_assign_stmt_472/type_cast_458_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_475/$entry
      -- CP-element group 124: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/$entry
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_1, ack => convTranspose_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	479 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Sample/ack
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_487_index_offset_ack_0, ack => convTranspose_CP_34_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	479 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_request/req
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_487_index_offset_ack_1, ack => convTranspose_CP_34_elements(126)); -- 
    req_995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(126), ack => addr_of_488_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_request/ack
      -- 
    ack_996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_488_final_reg_ack_0, ack => convTranspose_CP_34_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	479 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_complete/ack
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_488_final_reg_ack_1, ack => convTranspose_CP_34_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	479 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_update_start_
      -- CP-element group 129: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Update/cr
      -- 
    ra_1010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_491_inst_ack_0, ack => convTranspose_CP_34_elements(129)); -- 
    cr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(129), ack => RPIPE_ConvTranspose_input_pipe_491_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Sample/rr
      -- 
    ca_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_491_inst_ack_1, ack => convTranspose_CP_34_elements(130)); -- 
    rr_1023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => type_cast_495_inst_req_0); -- 
    rr_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => RPIPE_ConvTranspose_input_pipe_504_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Sample/ra
      -- 
    ra_1024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_495_inst_ack_0, ack => convTranspose_CP_34_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	479 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Update/ca
      -- 
    ca_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_495_inst_ack_1, ack => convTranspose_CP_34_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_update_start_
      -- CP-element group 133: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Update/cr
      -- 
    ra_1038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_504_inst_ack_0, ack => convTranspose_CP_34_elements(133)); -- 
    cr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(133), ack => RPIPE_ConvTranspose_input_pipe_504_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_504_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Sample/rr
      -- 
    ca_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_504_inst_ack_1, ack => convTranspose_CP_34_elements(134)); -- 
    rr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => type_cast_508_inst_req_0); -- 
    rr_1065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => RPIPE_ConvTranspose_input_pipe_522_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Sample/ra
      -- 
    ra_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_0, ack => convTranspose_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	479 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Update/ca
      -- 
    ca_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_1, ack => convTranspose_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_update_start_
      -- CP-element group 137: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Update/cr
      -- 
    ra_1066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_522_inst_ack_0, ack => convTranspose_CP_34_elements(137)); -- 
    cr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(137), ack => RPIPE_ConvTranspose_input_pipe_522_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_522_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Sample/rr
      -- 
    ca_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_522_inst_ack_1, ack => convTranspose_CP_34_elements(138)); -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => type_cast_526_inst_req_0); -- 
    rr_1093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => RPIPE_ConvTranspose_input_pipe_540_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Sample/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_526_inst_ack_0, ack => convTranspose_CP_34_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	479 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Update/ca
      -- 
    ca_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_526_inst_ack_1, ack => convTranspose_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_update_start_
      -- CP-element group 141: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_sample_completed_
      -- 
    ra_1094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_540_inst_ack_0, ack => convTranspose_CP_34_elements(141)); -- 
    cr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(141), ack => RPIPE_ConvTranspose_input_pipe_540_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_540_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Sample/$entry
      -- 
    ca_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_540_inst_ack_1, ack => convTranspose_CP_34_elements(142)); -- 
    rr_1107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => type_cast_544_inst_req_0); -- 
    rr_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => RPIPE_ConvTranspose_input_pipe_558_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_sample_completed_
      -- 
    ra_1108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_544_inst_ack_0, ack => convTranspose_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	479 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_update_completed_
      -- 
    ca_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_544_inst_ack_1, ack => convTranspose_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_update_start_
      -- CP-element group 145: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Sample/$exit
      -- 
    ra_1122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_558_inst_ack_0, ack => convTranspose_CP_34_elements(145)); -- 
    cr_1126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(145), ack => RPIPE_ConvTranspose_input_pipe_558_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_558_update_completed_
      -- 
    ca_1127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_558_inst_ack_1, ack => convTranspose_CP_34_elements(146)); -- 
    rr_1135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => type_cast_562_inst_req_0); -- 
    rr_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => RPIPE_ConvTranspose_input_pipe_576_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_sample_completed_
      -- 
    ra_1136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_562_inst_ack_0, ack => convTranspose_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	479 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_update_completed_
      -- 
    ca_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_562_inst_ack_1, ack => convTranspose_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_update_start_
      -- CP-element group 149: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_sample_completed_
      -- 
    ra_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_576_inst_ack_0, ack => convTranspose_CP_34_elements(149)); -- 
    cr_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(149), ack => RPIPE_ConvTranspose_input_pipe_576_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_576_update_completed_
      -- 
    ca_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_576_inst_ack_1, ack => convTranspose_CP_34_elements(150)); -- 
    rr_1163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => type_cast_580_inst_req_0); -- 
    rr_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => RPIPE_ConvTranspose_input_pipe_594_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_sample_completed_
      -- 
    ra_1164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_580_inst_ack_0, ack => convTranspose_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	479 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_update_completed_
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_580_inst_ack_1, ack => convTranspose_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_update_start_
      -- 
    ra_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_594_inst_ack_0, ack => convTranspose_CP_34_elements(153)); -- 
    cr_1182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(153), ack => RPIPE_ConvTranspose_input_pipe_594_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_594_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_sample_start_
      -- 
    ca_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_594_inst_ack_1, ack => convTranspose_CP_34_elements(154)); -- 
    rr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => type_cast_598_inst_req_0); -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => RPIPE_ConvTranspose_input_pipe_612_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_sample_completed_
      -- 
    ra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_0, ack => convTranspose_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	479 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Update/$exit
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_1, ack => convTranspose_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_update_start_
      -- CP-element group 157: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_sample_completed_
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_612_inst_ack_0, ack => convTranspose_CP_34_elements(157)); -- 
    cr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(157), ack => RPIPE_ConvTranspose_input_pipe_612_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_612_update_completed_
      -- 
    ca_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_612_inst_ack_1, ack => convTranspose_CP_34_elements(158)); -- 
    rr_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(158), ack => type_cast_616_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_sample_completed_
      -- 
    ra_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_0, ack => convTranspose_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	479 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_update_completed_
      -- 
    ca_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_1, ack => convTranspose_CP_34_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/ptr_deref_624_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/ptr_deref_624_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/ptr_deref_624_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/ptr_deref_624_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/$entry
      -- 
    rr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(161), ack => ptr_deref_624_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(128) & convTranspose_CP_34_elements(132) & convTranspose_CP_34_elements(136) & convTranspose_CP_34_elements(140) & convTranspose_CP_34_elements(144) & convTranspose_CP_34_elements(148) & convTranspose_CP_34_elements(152) & convTranspose_CP_34_elements(156) & convTranspose_CP_34_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_sample_completed_
      -- 
    ra_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_624_store_0_ack_0, ack => convTranspose_CP_34_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	479 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_update_completed_
      -- 
    ca_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_624_store_0_ack_1, ack => convTranspose_CP_34_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_39/R_exitcond3_639_place
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637__exit__
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638__entry__
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_39/if_stmt_638_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/$exit
      -- 
    branch_req_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(164), ack => if_stmt_638_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(163) & convTranspose_CP_34_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	473 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_39/if_stmt_638_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_39/merge_stmt_428__exit__
      -- CP-element group 165: 	 branch_block_stmt_39/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_39/if_stmt_638_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_39/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_39/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_39/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_39/merge_stmt_428_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_39/merge_stmt_428_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_39/merge_stmt_428_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_39/merge_stmt_428_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_39/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_39/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_638_branch_ack_1, ack => convTranspose_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	475 
    -- CP-element group 166: 	476 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_39/if_stmt_638_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_39/if_stmt_638_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_638_branch_ack_0, ack => convTranspose_CP_34_elements(166)); -- 
    rr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_481_inst_req_0); -- 
    cr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_481_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_sample_completed_
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_0, ack => convTranspose_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	480 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679__exit__
      -- CP-element group 168: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/type_cast_665_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_39/assign_stmt_650_to_assign_stmt_679/$exit
      -- CP-element group 168: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_682/$entry
      -- CP-element group 168: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/$entry
      -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_1, ack => convTranspose_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	485 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_sample_complete
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_694_index_offset_ack_0, ack => convTranspose_CP_34_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	485 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_request/req
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_base_plus_offset/$entry
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_694_index_offset_ack_1, ack => convTranspose_CP_34_elements(170)); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(170), ack => addr_of_695_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_request/ack
      -- CP-element group 171: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_request/$exit
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_695_final_reg_ack_0, ack => convTranspose_CP_34_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	485 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_word_addrgen/root_register_ack
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_695_final_reg_ack_1, ack => convTranspose_CP_34_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	485 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_update_start_
      -- CP-element group 173: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_sample_completed_
      -- 
    ra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_698_inst_ack_0, ack => convTranspose_CP_34_elements(173)); -- 
    cr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(173), ack => RPIPE_ConvTranspose_input_pipe_698_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Sample/$entry
      -- 
    ca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_698_inst_ack_1, ack => convTranspose_CP_34_elements(174)); -- 
    rr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => type_cast_702_inst_req_0); -- 
    rr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => RPIPE_ConvTranspose_input_pipe_711_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Sample/$exit
      -- 
    ra_1383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_702_inst_ack_0, ack => convTranspose_CP_34_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	485 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Update/$exit
      -- 
    ca_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_702_inst_ack_1, ack => convTranspose_CP_34_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_update_start_
      -- CP-element group 177: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_sample_completed_
      -- 
    ra_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_711_inst_ack_0, ack => convTranspose_CP_34_elements(177)); -- 
    cr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(177), ack => RPIPE_ConvTranspose_input_pipe_711_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_711_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Sample/$entry
      -- 
    ca_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_711_inst_ack_1, ack => convTranspose_CP_34_elements(178)); -- 
    rr_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => type_cast_715_inst_req_0); -- 
    rr_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => RPIPE_ConvTranspose_input_pipe_729_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Sample/$exit
      -- 
    ra_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_0, ack => convTranspose_CP_34_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	485 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Update/$exit
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_1, ack => convTranspose_CP_34_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_update_start_
      -- 
    ra_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_729_inst_ack_0, ack => convTranspose_CP_34_elements(181)); -- 
    cr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(181), ack => RPIPE_ConvTranspose_input_pipe_729_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_729_update_completed_
      -- 
    ca_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_729_inst_ack_1, ack => convTranspose_CP_34_elements(182)); -- 
    rr_1452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => RPIPE_ConvTranspose_input_pipe_747_inst_req_0); -- 
    rr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => type_cast_733_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Sample/ra
      -- 
    ra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_733_inst_ack_0, ack => convTranspose_CP_34_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	485 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Update/$exit
      -- 
    ca_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_733_inst_ack_1, ack => convTranspose_CP_34_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_update_start_
      -- 
    ra_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_747_inst_ack_0, ack => convTranspose_CP_34_elements(185)); -- 
    cr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(185), ack => RPIPE_ConvTranspose_input_pipe_747_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_747_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Sample/rr
      -- 
    ca_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_747_inst_ack_1, ack => convTranspose_CP_34_elements(186)); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => type_cast_751_inst_req_0); -- 
    rr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => RPIPE_ConvTranspose_input_pipe_765_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Sample/ra
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => convTranspose_CP_34_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	485 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Update/ca
      -- 
    ca_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => convTranspose_CP_34_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_update_start_
      -- CP-element group 189: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Update/cr
      -- 
    ra_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_765_inst_ack_0, ack => convTranspose_CP_34_elements(189)); -- 
    cr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(189), ack => RPIPE_ConvTranspose_input_pipe_765_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_765_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Sample/rr
      -- 
    ca_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_765_inst_ack_1, ack => convTranspose_CP_34_elements(190)); -- 
    rr_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => type_cast_769_inst_req_0); -- 
    rr_1508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => RPIPE_ConvTranspose_input_pipe_783_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Sample/ra
      -- 
    ra_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_0, ack => convTranspose_CP_34_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	485 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Update/ca
      -- 
    ca_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_1, ack => convTranspose_CP_34_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_update_start_
      -- CP-element group 193: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Update/cr
      -- 
    ra_1509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_783_inst_ack_0, ack => convTranspose_CP_34_elements(193)); -- 
    cr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(193), ack => RPIPE_ConvTranspose_input_pipe_783_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_783_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Sample/rr
      -- 
    ca_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_783_inst_ack_1, ack => convTranspose_CP_34_elements(194)); -- 
    rr_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => type_cast_787_inst_req_0); -- 
    rr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => RPIPE_ConvTranspose_input_pipe_801_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Sample/ra
      -- 
    ra_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_0, ack => convTranspose_CP_34_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	485 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Update/ca
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_1, ack => convTranspose_CP_34_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_update_start_
      -- CP-element group 197: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Update/cr
      -- 
    ra_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_801_inst_ack_0, ack => convTranspose_CP_34_elements(197)); -- 
    cr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(197), ack => RPIPE_ConvTranspose_input_pipe_801_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_801_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Sample/rr
      -- 
    ca_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_801_inst_ack_1, ack => convTranspose_CP_34_elements(198)); -- 
    rr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => type_cast_805_inst_req_0); -- 
    rr_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => RPIPE_ConvTranspose_input_pipe_819_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Sample/ra
      -- 
    ra_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_805_inst_ack_0, ack => convTranspose_CP_34_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	485 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Update/ca
      -- 
    ca_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_805_inst_ack_1, ack => convTranspose_CP_34_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_update_start_
      -- CP-element group 201: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Update/cr
      -- 
    ra_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_819_inst_ack_0, ack => convTranspose_CP_34_elements(201)); -- 
    cr_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(201), ack => RPIPE_ConvTranspose_input_pipe_819_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_819_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Sample/rr
      -- 
    ca_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_819_inst_ack_1, ack => convTranspose_CP_34_elements(202)); -- 
    rr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(202), ack => type_cast_823_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Sample/ra
      -- 
    ra_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_0, ack => convTranspose_CP_34_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	485 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Update/ca
      -- 
    ca_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_1, ack => convTranspose_CP_34_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/ptr_deref_831_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/ptr_deref_831_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/ptr_deref_831_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/ptr_deref_831_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/word_access_start/word_0/rr
      -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(205), ack => ptr_deref_831_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(184) & convTranspose_CP_34_elements(188) & convTranspose_CP_34_elements(192) & convTranspose_CP_34_elements(196) & convTranspose_CP_34_elements(200) & convTranspose_CP_34_elements(204) & convTranspose_CP_34_elements(180) & convTranspose_CP_34_elements(172) & convTranspose_CP_34_elements(176);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Sample/word_access_start/word_0/ra
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_831_store_0_ack_0, ack => convTranspose_CP_34_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	485 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/word_access_complete/word_0/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_831_store_0_ack_1, ack => convTranspose_CP_34_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844__exit__
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845__entry__
      -- CP-element group 208: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/$exit
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_39/R_exitcond2_846_place
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_39/if_stmt_845_else_link/$entry
      -- 
    branch_req_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(208), ack => if_stmt_845_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(207) & convTranspose_CP_34_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	486 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_39/merge_stmt_851__exit__
      -- CP-element group 209: 	 branch_block_stmt_39/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_39/if_stmt_845_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_39/if_stmt_845_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_39/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_39/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_39/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_39/merge_stmt_851_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_39/merge_stmt_851_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_39/merge_stmt_851_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_39/merge_stmt_851_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_39/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_39/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_845_branch_ack_1, ack => convTranspose_CP_34_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	481 
    -- CP-element group 210: 	482 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_39/if_stmt_845_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_39/if_stmt_845_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_845_branch_ack_0, ack => convTranspose_CP_34_elements(210)); -- 
    rr_3579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_685_inst_req_0); -- 
    cr_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_685_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	486 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Sample/ra
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_856_inst_ack_0, ack => convTranspose_CP_34_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	486 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Update/ca
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_856_inst_ack_1, ack => convTranspose_CP_34_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	486 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_0, ack => convTranspose_CP_34_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	486 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_1, ack => convTranspose_CP_34_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	486 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_864_inst_ack_0, ack => convTranspose_CP_34_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	486 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_864_inst_ack_1, ack => convTranspose_CP_34_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881__exit__
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882__entry__
      -- CP-element group 217: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/$exit
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_39/R_cmp264506_883_place
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_39/if_stmt_882_else_link/$entry
      -- 
    branch_req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(217), ack => if_stmt_882_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(212) & convTranspose_CP_34_elements(214) & convTranspose_CP_34_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_39/merge_stmt_888__exit__
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923__entry__
      -- CP-element group 218: 	 branch_block_stmt_39/if_stmt_882_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_39/if_stmt_882_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_39/forx_xend250_bbx_xnph508
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/$entry
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_update_start_
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_39/forx_xend250_bbx_xnph508_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_39/forx_xend250_bbx_xnph508_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_39/merge_stmt_888_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_39/merge_stmt_888_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_39/merge_stmt_888_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_39/merge_stmt_888_PhiAck/dummy
      -- 
    if_choice_transition_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_882_branch_ack_1, ack => convTranspose_CP_34_elements(218)); -- 
    rr_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_909_inst_req_0); -- 
    cr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_909_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	493 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_39/if_stmt_882_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_39/if_stmt_882_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_39/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_39/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_39/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_882_branch_ack_0, ack => convTranspose_CP_34_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Sample/ra
      -- 
    ra_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_909_inst_ack_0, ack => convTranspose_CP_34_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	487 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923__exit__
      -- CP-element group 221: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/$exit
      -- CP-element group 221: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_39/assign_stmt_894_to_assign_stmt_923/type_cast_909_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_926/$entry
      -- CP-element group 221: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/$entry
      -- 
    ca_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_909_inst_ack_1, ack => convTranspose_CP_34_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	492 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Sample/ack
      -- 
    ack_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_offset_ack_0, ack => convTranspose_CP_34_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	492 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_request/req
      -- 
    ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_offset_ack_1, ack => convTranspose_CP_34_elements(223)); -- 
    req_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(223), ack => addr_of_939_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_request/ack
      -- 
    ack_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_939_final_reg_ack_0, ack => convTranspose_CP_34_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	492 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/ptr_deref_942_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/ptr_deref_942_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/ptr_deref_942_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/ptr_deref_942_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/word_access_start/word_0/rr
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_939_final_reg_ack_1, ack => convTranspose_CP_34_elements(225)); -- 
    rr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(225), ack => ptr_deref_942_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Sample/word_access_start/word_0/ra
      -- 
    ra_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_942_store_0_ack_0, ack => convTranspose_CP_34_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	492 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/word_access_complete/word_0/ca
      -- 
    ca_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_942_store_0_ack_1, ack => convTranspose_CP_34_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956__exit__
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957__entry__
      -- CP-element group 228: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/$exit
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_39/R_exitcond_958_place
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_39/if_stmt_957_else_link/$entry
      -- 
    branch_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(228), ack => if_stmt_957_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(222) & convTranspose_CP_34_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	493 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_39/merge_stmt_963__exit__
      -- CP-element group 229: 	 branch_block_stmt_39/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_39/if_stmt_957_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_39/if_stmt_957_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_39/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_39/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_39/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_39/merge_stmt_963_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_39/merge_stmt_963_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_39/merge_stmt_963_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_39/merge_stmt_963_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_39/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_39/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_957_branch_ack_1, ack => convTranspose_CP_34_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	488 
    -- CP-element group 230: 	489 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_39/if_stmt_957_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_39/if_stmt_957_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_957_branch_ack_0, ack => convTranspose_CP_34_elements(230)); -- 
    rr_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_929_inst_req_0); -- 
    cr_3661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_929_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	493 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Sample/cra
      -- 
    cra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_968_call_ack_0, ack => convTranspose_CP_34_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	493 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Sample/rr
      -- 
    cca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_968_call_ack_1, ack => convTranspose_CP_34_elements(232)); -- 
    rr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(232), ack => type_cast_973_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Sample/ra
      -- 
    ra_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_973_inst_ack_0, ack => convTranspose_CP_34_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	493 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	349 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234:  members (55) 
      -- CP-element group 234: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974__exit__
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187__entry__
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_update_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_update_start_
      -- CP-element group 234: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/$exit
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_update_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_update_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_update_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_update_start_
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Update/cr
      -- 
    ca_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_973_inst_ack_1, ack => convTranspose_CP_34_elements(234)); -- 
    req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block2_start_1076_inst_req_0); -- 
    rr_2216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1055_inst_req_0); -- 
    cr_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1055_inst_req_1); -- 
    req_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block1_start_1020_inst_req_0); -- 
    cr_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1062_inst_req_1); -- 
    rr_2244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1062_inst_req_0); -- 
    req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block0_start_976_inst_req_0); -- 
    rr_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1111_inst_req_0); -- 
    cr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1111_inst_req_1); -- 
    rr_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1118_inst_req_0); -- 
    cr_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1118_inst_req_1); -- 
    req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block3_start_1132_inst_req_0); -- 
    rr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1167_inst_req_0); -- 
    cr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1167_inst_req_1); -- 
    rr_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1174_inst_req_0); -- 
    cr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1174_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_update_start_
      -- CP-element group 235: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Update/req
      -- 
    ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_0, ack => convTranspose_CP_34_elements(235)); -- 
    req_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(235), ack => WPIPE_Block0_start_976_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_976_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_sample_start_
      -- 
    ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_1, ack => convTranspose_CP_34_elements(236)); -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(236), ack => WPIPE_Block0_start_979_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Update/req
      -- CP-element group 237: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_update_start_
      -- CP-element group 237: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_sample_completed_
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_0, ack => convTranspose_CP_34_elements(237)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(237), ack => WPIPE_Block0_start_979_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_979_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Sample/req
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_1, ack => convTranspose_CP_34_elements(238)); -- 
    req_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(238), ack => WPIPE_Block0_start_982_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_update_start_
      -- CP-element group 239: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Update/req
      -- CP-element group 239: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Sample/ack
      -- 
    ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_0, ack => convTranspose_CP_34_elements(239)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(239), ack => WPIPE_Block0_start_982_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Sample/req
      -- CP-element group 240: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_982_Update/$exit
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_1, ack => convTranspose_CP_34_elements(240)); -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(240), ack => WPIPE_Block0_start_985_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Update/req
      -- CP-element group 241: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_update_start_
      -- CP-element group 241: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_sample_completed_
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_0, ack => convTranspose_CP_34_elements(241)); -- 
    req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(241), ack => WPIPE_Block0_start_985_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_985_update_completed_
      -- 
    ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_1, ack => convTranspose_CP_34_elements(242)); -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(242), ack => WPIPE_Block0_start_988_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_update_start_
      -- CP-element group 243: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Update/req
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_0, ack => convTranspose_CP_34_elements(243)); -- 
    req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(243), ack => WPIPE_Block0_start_988_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_988_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Sample/req
      -- 
    ack_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_1, ack => convTranspose_CP_34_elements(244)); -- 
    req_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(244), ack => WPIPE_Block0_start_991_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_update_start_
      -- CP-element group 245: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Update/req
      -- CP-element group 245: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Sample/ack
      -- 
    ack_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_991_inst_ack_0, ack => convTranspose_CP_34_elements(245)); -- 
    req_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(245), ack => WPIPE_Block0_start_991_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_991_Update/$exit
      -- 
    ack_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_991_inst_ack_1, ack => convTranspose_CP_34_elements(246)); -- 
    req_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(246), ack => WPIPE_Block0_start_994_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Update/req
      -- CP-element group 247: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_update_start_
      -- CP-element group 247: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_sample_completed_
      -- 
    ack_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_0, ack => convTranspose_CP_34_elements(247)); -- 
    req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(247), ack => WPIPE_Block0_start_994_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_994_update_completed_
      -- 
    ack_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_1, ack => convTranspose_CP_34_elements(248)); -- 
    req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(248), ack => WPIPE_Block0_start_997_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_update_start_
      -- CP-element group 249: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Update/req
      -- 
    ack_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_997_inst_ack_0, ack => convTranspose_CP_34_elements(249)); -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(249), ack => WPIPE_Block0_start_997_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_997_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Sample/req
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_997_inst_ack_1, ack => convTranspose_CP_34_elements(250)); -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(250), ack => WPIPE_Block0_start_1000_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_update_start_
      -- CP-element group 251: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Update/req
      -- CP-element group 251: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Update/$entry
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1000_inst_ack_0, ack => convTranspose_CP_34_elements(251)); -- 
    req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(251), ack => WPIPE_Block0_start_1000_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1000_Update/$exit
      -- 
    ack_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1000_inst_ack_1, ack => convTranspose_CP_34_elements(252)); -- 
    req_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(252), ack => WPIPE_Block0_start_1003_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Update/req
      -- CP-element group 253: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_update_start_
      -- CP-element group 253: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_sample_completed_
      -- 
    ack_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1003_inst_ack_0, ack => convTranspose_CP_34_elements(253)); -- 
    req_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(253), ack => WPIPE_Block0_start_1003_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1003_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Sample/$entry
      -- 
    ack_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1003_inst_ack_1, ack => convTranspose_CP_34_elements(254)); -- 
    req_2034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(254), ack => WPIPE_Block0_start_1007_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_update_start_
      -- CP-element group 255: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Update/req
      -- CP-element group 255: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Sample/$exit
      -- 
    ack_2035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1007_inst_ack_0, ack => convTranspose_CP_34_elements(255)); -- 
    req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(255), ack => WPIPE_Block0_start_1007_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1007_update_completed_
      -- 
    ack_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1007_inst_ack_1, ack => convTranspose_CP_34_elements(256)); -- 
    req_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(256), ack => WPIPE_Block0_start_1011_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Update/req
      -- CP-element group 257: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_update_start_
      -- CP-element group 257: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_sample_completed_
      -- 
    ack_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1011_inst_ack_0, ack => convTranspose_CP_34_elements(257)); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(257), ack => WPIPE_Block0_start_1011_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1011_update_completed_
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1011_inst_ack_1, ack => convTranspose_CP_34_elements(258)); -- 
    req_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(258), ack => WPIPE_Block0_start_1014_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Update/req
      -- CP-element group 259: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_update_start_
      -- CP-element group 259: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_sample_completed_
      -- 
    ack_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1014_inst_ack_0, ack => convTranspose_CP_34_elements(259)); -- 
    req_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(259), ack => WPIPE_Block0_start_1014_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1014_update_completed_
      -- 
    ack_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1014_inst_ack_1, ack => convTranspose_CP_34_elements(260)); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(260), ack => WPIPE_Block0_start_1017_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Update/req
      -- CP-element group 261: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_update_start_
      -- CP-element group 261: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_sample_completed_
      -- 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1017_inst_ack_0, ack => convTranspose_CP_34_elements(261)); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(261), ack => WPIPE_Block0_start_1017_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	365 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block0_start_1017_Update/ack
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1017_inst_ack_1, ack => convTranspose_CP_34_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_update_start_
      -- CP-element group 263: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Update/req
      -- 
    ack_2091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1020_inst_ack_0, ack => convTranspose_CP_34_elements(263)); -- 
    req_2095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(263), ack => WPIPE_Block1_start_1020_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1020_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Sample/req
      -- 
    ack_2096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1020_inst_ack_1, ack => convTranspose_CP_34_elements(264)); -- 
    req_2104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => WPIPE_Block1_start_1023_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_update_start_
      -- CP-element group 265: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Update/req
      -- 
    ack_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1023_inst_ack_0, ack => convTranspose_CP_34_elements(265)); -- 
    req_2109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(265), ack => WPIPE_Block1_start_1023_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1023_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Sample/$entry
      -- 
    ack_2110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1023_inst_ack_1, ack => convTranspose_CP_34_elements(266)); -- 
    req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(266), ack => WPIPE_Block1_start_1026_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Update/req
      -- CP-element group 267: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_update_start_
      -- CP-element group 267: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_sample_completed_
      -- 
    ack_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1026_inst_ack_0, ack => convTranspose_CP_34_elements(267)); -- 
    req_2123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(267), ack => WPIPE_Block1_start_1026_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1026_update_completed_
      -- 
    ack_2124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1026_inst_ack_1, ack => convTranspose_CP_34_elements(268)); -- 
    req_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => WPIPE_Block1_start_1029_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Update/req
      -- CP-element group 269: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_update_start_
      -- CP-element group 269: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_sample_completed_
      -- 
    ack_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1029_inst_ack_0, ack => convTranspose_CP_34_elements(269)); -- 
    req_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(269), ack => WPIPE_Block1_start_1029_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1029_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Sample/req
      -- 
    ack_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1029_inst_ack_1, ack => convTranspose_CP_34_elements(270)); -- 
    req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(270), ack => WPIPE_Block1_start_1032_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_update_start_
      -- CP-element group 271: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Update/req
      -- CP-element group 271: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Sample/ack
      -- 
    ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1032_inst_ack_0, ack => convTranspose_CP_34_elements(271)); -- 
    req_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(271), ack => WPIPE_Block1_start_1032_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1032_Update/$exit
      -- 
    ack_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1032_inst_ack_1, ack => convTranspose_CP_34_elements(272)); -- 
    req_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(272), ack => WPIPE_Block1_start_1035_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Update/req
      -- CP-element group 273: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_update_start_
      -- CP-element group 273: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_sample_completed_
      -- 
    ack_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1035_inst_ack_0, ack => convTranspose_CP_34_elements(273)); -- 
    req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(273), ack => WPIPE_Block1_start_1035_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1035_update_completed_
      -- 
    ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1035_inst_ack_1, ack => convTranspose_CP_34_elements(274)); -- 
    req_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(274), ack => WPIPE_Block1_start_1038_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Update/req
      -- CP-element group 275: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_update_start_
      -- CP-element group 275: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_sample_completed_
      -- 
    ack_2175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1038_inst_ack_0, ack => convTranspose_CP_34_elements(275)); -- 
    req_2179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(275), ack => WPIPE_Block1_start_1038_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1038_update_completed_
      -- 
    ack_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1038_inst_ack_1, ack => convTranspose_CP_34_elements(276)); -- 
    req_2188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(276), ack => WPIPE_Block1_start_1041_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Update/req
      -- CP-element group 277: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_update_start_
      -- CP-element group 277: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_sample_completed_
      -- 
    ack_2189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1041_inst_ack_0, ack => convTranspose_CP_34_elements(277)); -- 
    req_2193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(277), ack => WPIPE_Block1_start_1041_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1041_update_completed_
      -- 
    ack_2194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1041_inst_ack_1, ack => convTranspose_CP_34_elements(278)); -- 
    req_2202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(278), ack => WPIPE_Block1_start_1044_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_update_start_
      -- CP-element group 279: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Update/req
      -- CP-element group 279: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_sample_completed_
      -- 
    ack_2203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1044_inst_ack_0, ack => convTranspose_CP_34_elements(279)); -- 
    req_2207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(279), ack => WPIPE_Block1_start_1044_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1044_Update/$exit
      -- 
    ack_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1044_inst_ack_1, ack => convTranspose_CP_34_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Sample/ra
      -- 
    ra_2217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => convTranspose_CP_34_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1055_Update/ca
      -- 
    ca_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => convTranspose_CP_34_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Sample/req
      -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(283), ack => WPIPE_Block1_start_1057_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(280) & convTranspose_CP_34_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Update/req
      -- CP-element group 284: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_update_start_
      -- CP-element group 284: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Update/$entry
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_0, ack => convTranspose_CP_34_elements(284)); -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(284), ack => WPIPE_Block1_start_1057_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1057_Update/ack
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_1, ack => convTranspose_CP_34_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_sample_completed_
      -- 
    ra_2245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_0, ack => convTranspose_CP_34_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1062_update_completed_
      -- 
    ca_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_1, ack => convTranspose_CP_34_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_sample_start_
      -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(288), ack => WPIPE_Block1_start_1064_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(285) & convTranspose_CP_34_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Update/req
      -- CP-element group 289: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_update_start_
      -- CP-element group 289: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_sample_completed_
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1064_inst_ack_0, ack => convTranspose_CP_34_elements(289)); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(289), ack => WPIPE_Block1_start_1064_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1064_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Sample/$entry
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1064_inst_ack_1, ack => convTranspose_CP_34_elements(290)); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(290), ack => WPIPE_Block1_start_1067_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Update/req
      -- CP-element group 291: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_update_start_
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1067_inst_ack_0, ack => convTranspose_CP_34_elements(291)); -- 
    req_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(291), ack => WPIPE_Block1_start_1067_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1067_update_completed_
      -- 
    ack_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1067_inst_ack_1, ack => convTranspose_CP_34_elements(292)); -- 
    req_2286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(292), ack => WPIPE_Block1_start_1070_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Update/req
      -- CP-element group 293: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_update_start_
      -- CP-element group 293: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Sample/$exit
      -- 
    ack_2287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1070_inst_ack_0, ack => convTranspose_CP_34_elements(293)); -- 
    req_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(293), ack => WPIPE_Block1_start_1070_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1070_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_sample_start_
      -- 
    ack_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1070_inst_ack_1, ack => convTranspose_CP_34_elements(294)); -- 
    req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(294), ack => WPIPE_Block1_start_1073_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Update/req
      -- CP-element group 295: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_update_start_
      -- CP-element group 295: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_sample_completed_
      -- 
    ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1073_inst_ack_0, ack => convTranspose_CP_34_elements(295)); -- 
    req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(295), ack => WPIPE_Block1_start_1073_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	365 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block1_start_1073_update_completed_
      -- 
    ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1073_inst_ack_1, ack => convTranspose_CP_34_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_update_start_
      -- CP-element group 297: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Update/req
      -- CP-element group 297: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Update/$entry
      -- 
    ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1076_inst_ack_0, ack => convTranspose_CP_34_elements(297)); -- 
    req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(297), ack => WPIPE_Block2_start_1076_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1076_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Sample/$entry
      -- 
    ack_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1076_inst_ack_1, ack => convTranspose_CP_34_elements(298)); -- 
    req_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(298), ack => WPIPE_Block2_start_1079_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_update_start_
      -- CP-element group 299: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Update/req
      -- CP-element group 299: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Sample/$exit
      -- 
    ack_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1079_inst_ack_0, ack => convTranspose_CP_34_elements(299)); -- 
    req_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(299), ack => WPIPE_Block2_start_1079_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1079_update_completed_
      -- 
    ack_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1079_inst_ack_1, ack => convTranspose_CP_34_elements(300)); -- 
    req_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(300), ack => WPIPE_Block2_start_1082_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_update_start_
      -- CP-element group 301: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Update/req
      -- CP-element group 301: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Sample/$exit
      -- 
    ack_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1082_inst_ack_0, ack => convTranspose_CP_34_elements(301)); -- 
    req_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(301), ack => WPIPE_Block2_start_1082_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1082_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_sample_start_
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1082_inst_ack_1, ack => convTranspose_CP_34_elements(302)); -- 
    req_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(302), ack => WPIPE_Block2_start_1085_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Update/req
      -- CP-element group 303: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_update_start_
      -- CP-element group 303: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_sample_completed_
      -- 
    ack_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1085_inst_ack_0, ack => convTranspose_CP_34_elements(303)); -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(303), ack => WPIPE_Block2_start_1085_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1085_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Sample/$entry
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1085_inst_ack_1, ack => convTranspose_CP_34_elements(304)); -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(304), ack => WPIPE_Block2_start_1088_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Update/req
      -- CP-element group 305: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_update_start_
      -- CP-element group 305: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Sample/$exit
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1088_inst_ack_0, ack => convTranspose_CP_34_elements(305)); -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(305), ack => WPIPE_Block2_start_1088_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1088_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_sample_start_
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1088_inst_ack_1, ack => convTranspose_CP_34_elements(306)); -- 
    req_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(306), ack => WPIPE_Block2_start_1091_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_update_start_
      -- CP-element group 307: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Update/req
      -- CP-element group 307: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Update/$entry
      -- 
    ack_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1091_inst_ack_0, ack => convTranspose_CP_34_elements(307)); -- 
    req_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(307), ack => WPIPE_Block2_start_1091_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1091_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Sample/req
      -- 
    ack_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1091_inst_ack_1, ack => convTranspose_CP_34_elements(308)); -- 
    req_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(308), ack => WPIPE_Block2_start_1094_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_update_start_
      -- CP-element group 309: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Update/req
      -- 
    ack_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1094_inst_ack_0, ack => convTranspose_CP_34_elements(309)); -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(309), ack => WPIPE_Block2_start_1094_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1094_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Sample/req
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1094_inst_ack_1, ack => convTranspose_CP_34_elements(310)); -- 
    req_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(310), ack => WPIPE_Block2_start_1097_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_update_start_
      -- CP-element group 311: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Update/req
      -- 
    ack_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1097_inst_ack_0, ack => convTranspose_CP_34_elements(311)); -- 
    req_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(311), ack => WPIPE_Block2_start_1097_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1097_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Sample/req
      -- 
    ack_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1097_inst_ack_1, ack => convTranspose_CP_34_elements(312)); -- 
    req_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(312), ack => WPIPE_Block2_start_1100_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_update_start_
      -- CP-element group 313: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Update/req
      -- 
    ack_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1100_inst_ack_0, ack => convTranspose_CP_34_elements(313)); -- 
    req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(313), ack => WPIPE_Block2_start_1100_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1100_Update/ack
      -- 
    ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1100_inst_ack_1, ack => convTranspose_CP_34_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Sample/ra
      -- 
    ra_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_0, ack => convTranspose_CP_34_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1111_Update/ca
      -- 
    ca_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_1, ack => convTranspose_CP_34_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Sample/req
      -- 
    req_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => WPIPE_Block2_start_1113_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(314) & convTranspose_CP_34_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_update_start_
      -- CP-element group 318: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Update/req
      -- 
    ack_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_0, ack => convTranspose_CP_34_elements(318)); -- 
    req_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(318), ack => WPIPE_Block2_start_1113_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1113_Update/ack
      -- 
    ack_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_1, ack => convTranspose_CP_34_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Sample/ra
      -- 
    ra_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1118_inst_ack_0, ack => convTranspose_CP_34_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1118_Update/ca
      -- 
    ca_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1118_inst_ack_1, ack => convTranspose_CP_34_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Sample/req
      -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(322), ack => WPIPE_Block2_start_1120_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(319) & convTranspose_CP_34_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_update_start_
      -- CP-element group 323: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Update/req
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1120_inst_ack_0, ack => convTranspose_CP_34_elements(323)); -- 
    req_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(323), ack => WPIPE_Block2_start_1120_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1120_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Sample/req
      -- 
    ack_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1120_inst_ack_1, ack => convTranspose_CP_34_elements(324)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(324), ack => WPIPE_Block2_start_1123_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_update_start_
      -- CP-element group 325: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Update/req
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1123_inst_ack_0, ack => convTranspose_CP_34_elements(325)); -- 
    req_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(325), ack => WPIPE_Block2_start_1123_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1123_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Sample/req
      -- 
    ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1123_inst_ack_1, ack => convTranspose_CP_34_elements(326)); -- 
    req_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(326), ack => WPIPE_Block2_start_1126_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_update_start_
      -- CP-element group 327: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Update/req
      -- 
    ack_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1126_inst_ack_0, ack => convTranspose_CP_34_elements(327)); -- 
    req_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(327), ack => WPIPE_Block2_start_1126_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1126_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Sample/req
      -- 
    ack_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1126_inst_ack_1, ack => convTranspose_CP_34_elements(328)); -- 
    req_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(328), ack => WPIPE_Block2_start_1129_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_update_start_
      -- CP-element group 329: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Update/req
      -- 
    ack_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1129_inst_ack_0, ack => convTranspose_CP_34_elements(329)); -- 
    req_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(329), ack => WPIPE_Block2_start_1129_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	365 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block2_start_1129_Update/ack
      -- 
    ack_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1129_inst_ack_1, ack => convTranspose_CP_34_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_update_start_
      -- CP-element group 331: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Update/req
      -- 
    ack_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1132_inst_ack_0, ack => convTranspose_CP_34_elements(331)); -- 
    req_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(331), ack => WPIPE_Block3_start_1132_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1132_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Sample/req
      -- 
    ack_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1132_inst_ack_1, ack => convTranspose_CP_34_elements(332)); -- 
    req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(332), ack => WPIPE_Block3_start_1135_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_update_start_
      -- CP-element group 333: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Update/req
      -- 
    ack_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1135_inst_ack_0, ack => convTranspose_CP_34_elements(333)); -- 
    req_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(333), ack => WPIPE_Block3_start_1135_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1135_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Sample/req
      -- 
    ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1135_inst_ack_1, ack => convTranspose_CP_34_elements(334)); -- 
    req_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(334), ack => WPIPE_Block3_start_1138_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_update_start_
      -- CP-element group 335: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Update/req
      -- 
    ack_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1138_inst_ack_0, ack => convTranspose_CP_34_elements(335)); -- 
    req_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(335), ack => WPIPE_Block3_start_1138_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1138_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Sample/req
      -- 
    ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1138_inst_ack_1, ack => convTranspose_CP_34_elements(336)); -- 
    req_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(336), ack => WPIPE_Block3_start_1141_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_update_start_
      -- CP-element group 337: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Update/req
      -- 
    ack_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1141_inst_ack_0, ack => convTranspose_CP_34_elements(337)); -- 
    req_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(337), ack => WPIPE_Block3_start_1141_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1141_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Sample/req
      -- 
    ack_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1141_inst_ack_1, ack => convTranspose_CP_34_elements(338)); -- 
    req_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(338), ack => WPIPE_Block3_start_1144_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_update_start_
      -- CP-element group 339: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Update/req
      -- 
    ack_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1144_inst_ack_0, ack => convTranspose_CP_34_elements(339)); -- 
    req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(339), ack => WPIPE_Block3_start_1144_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1144_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Sample/req
      -- 
    ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1144_inst_ack_1, ack => convTranspose_CP_34_elements(340)); -- 
    req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(340), ack => WPIPE_Block3_start_1147_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_update_start_
      -- CP-element group 341: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Update/req
      -- 
    ack_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1147_inst_ack_0, ack => convTranspose_CP_34_elements(341)); -- 
    req_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(341), ack => WPIPE_Block3_start_1147_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1147_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Sample/req
      -- 
    ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1147_inst_ack_1, ack => convTranspose_CP_34_elements(342)); -- 
    req_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(342), ack => WPIPE_Block3_start_1150_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_update_start_
      -- CP-element group 343: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Update/req
      -- 
    ack_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1150_inst_ack_0, ack => convTranspose_CP_34_elements(343)); -- 
    req_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(343), ack => WPIPE_Block3_start_1150_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1150_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Sample/req
      -- 
    ack_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1150_inst_ack_1, ack => convTranspose_CP_34_elements(344)); -- 
    req_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(344), ack => WPIPE_Block3_start_1153_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_update_start_
      -- CP-element group 345: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Update/req
      -- 
    ack_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1153_inst_ack_0, ack => convTranspose_CP_34_elements(345)); -- 
    req_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(345), ack => WPIPE_Block3_start_1153_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1153_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Sample/req
      -- 
    ack_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1153_inst_ack_1, ack => convTranspose_CP_34_elements(346)); -- 
    req_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(346), ack => WPIPE_Block3_start_1156_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_update_start_
      -- CP-element group 347: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Update/req
      -- 
    ack_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1156_inst_ack_0, ack => convTranspose_CP_34_elements(347)); -- 
    req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(347), ack => WPIPE_Block3_start_1156_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1156_Update/ack
      -- 
    ack_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1156_inst_ack_1, ack => convTranspose_CP_34_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Sample/ra
      -- 
    ra_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => convTranspose_CP_34_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1167_Update/ca
      -- 
    ca_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => convTranspose_CP_34_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Sample/req
      -- 
    req_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(351), ack => WPIPE_Block3_start_1169_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(348) & convTranspose_CP_34_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_update_start_
      -- CP-element group 352: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Update/req
      -- 
    ack_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_0, ack => convTranspose_CP_34_elements(352)); -- 
    req_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(352), ack => WPIPE_Block3_start_1169_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1169_Update/ack
      -- 
    ack_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_1, ack => convTranspose_CP_34_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Sample/ra
      -- 
    ra_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_0, ack => convTranspose_CP_34_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/type_cast_1174_Update/ca
      -- 
    ca_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_1, ack => convTranspose_CP_34_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Sample/req
      -- 
    req_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(356), ack => WPIPE_Block3_start_1176_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(353) & convTranspose_CP_34_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_update_start_
      -- CP-element group 357: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Update/req
      -- 
    ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1176_inst_ack_0, ack => convTranspose_CP_34_elements(357)); -- 
    req_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(357), ack => WPIPE_Block3_start_1176_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1176_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Sample/req
      -- 
    ack_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1176_inst_ack_1, ack => convTranspose_CP_34_elements(358)); -- 
    req_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(358), ack => WPIPE_Block3_start_1179_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_update_start_
      -- CP-element group 359: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Update/req
      -- 
    ack_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1179_inst_ack_0, ack => convTranspose_CP_34_elements(359)); -- 
    req_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(359), ack => WPIPE_Block3_start_1179_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1179_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Sample/req
      -- 
    ack_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1179_inst_ack_1, ack => convTranspose_CP_34_elements(360)); -- 
    req_2734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(360), ack => WPIPE_Block3_start_1182_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_update_start_
      -- CP-element group 361: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Update/req
      -- 
    ack_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1182_inst_ack_0, ack => convTranspose_CP_34_elements(361)); -- 
    req_2739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(361), ack => WPIPE_Block3_start_1182_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1182_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Sample/req
      -- 
    ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1182_inst_ack_1, ack => convTranspose_CP_34_elements(362)); -- 
    req_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(362), ack => WPIPE_Block3_start_1185_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_update_start_
      -- CP-element group 363: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Update/req
      -- 
    ack_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1185_inst_ack_0, ack => convTranspose_CP_34_elements(363)); -- 
    req_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(363), ack => WPIPE_Block3_start_1185_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/WPIPE_Block3_start_1185_Update/ack
      -- 
    ack_2754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1185_inst_ack_1, ack => convTranspose_CP_34_elements(364)); -- 
    -- CP-element group 365:  join  fork  transition  place  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	262 
    -- CP-element group 365: 	296 
    -- CP-element group 365: 	330 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: 	368 
    -- CP-element group 365: 	370 
    -- CP-element group 365: 	372 
    -- CP-element group 365:  members (16) 
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187__exit__
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200__entry__
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_978_to_assign_stmt_1187/$exit
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/$entry
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Sample/rr
      -- 
    rr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block0_done_1190_inst_req_0); -- 
    rr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block1_done_1193_inst_req_0); -- 
    rr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block2_done_1196_inst_req_0); -- 
    rr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block3_done_1199_inst_req_0); -- 
    convTranspose_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(262) & convTranspose_CP_34_elements(296) & convTranspose_CP_34_elements(330) & convTranspose_CP_34_elements(364);
      gj_convTranspose_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (6) 
      -- CP-element group 366: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_update_start_
      -- CP-element group 366: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Sample/ra
      -- CP-element group 366: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Update/cr
      -- 
    ra_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1190_inst_ack_0, ack => convTranspose_CP_34_elements(366)); -- 
    cr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => RPIPE_Block0_done_1190_inst_req_1); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	374 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block0_done_1190_Update/ca
      -- 
    ca_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1190_inst_ack_1, ack => convTranspose_CP_34_elements(367)); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	365 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_update_start_
      -- CP-element group 368: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Sample/ra
      -- CP-element group 368: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Update/cr
      -- 
    ra_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1193_inst_ack_0, ack => convTranspose_CP_34_elements(368)); -- 
    cr_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(368), ack => RPIPE_Block1_done_1193_inst_req_1); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block1_done_1193_Update/ca
      -- 
    ca_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1193_inst_ack_1, ack => convTranspose_CP_34_elements(369)); -- 
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_update_start_
      -- CP-element group 370: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Sample/ra
      -- CP-element group 370: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Update/cr
      -- 
    ra_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1196_inst_ack_0, ack => convTranspose_CP_34_elements(370)); -- 
    cr_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(370), ack => RPIPE_Block2_done_1196_inst_req_1); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	374 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block2_done_1196_Update/ca
      -- 
    ca_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1196_inst_ack_1, ack => convTranspose_CP_34_elements(371)); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	365 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_update_start_
      -- CP-element group 372: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Sample/ra
      -- CP-element group 372: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Update/cr
      -- 
    ra_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1199_inst_ack_0, ack => convTranspose_CP_34_elements(372)); -- 
    cr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => RPIPE_Block3_done_1199_inst_req_1); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/RPIPE_Block3_done_1199_Update/ca
      -- 
    ca_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1199_inst_ack_1, ack => convTranspose_CP_34_elements(373)); -- 
    -- CP-element group 374:  join  fork  transition  place  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	367 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	371 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	384 
    -- CP-element group 374: 	386 
    -- CP-element group 374: 	388 
    -- CP-element group 374: 	390 
    -- CP-element group 374: 	392 
    -- CP-element group 374: 	394 
    -- CP-element group 374: 	396 
    -- CP-element group 374: 	378 
    -- CP-element group 374: 	382 
    -- CP-element group 374: 	375 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (37) 
      -- CP-element group 374: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200__exit__
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314__entry__
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/assign_stmt_1191_to_assign_stmt_1200/$exit
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Sample/crr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Update/ccr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_update_start_
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_update_start_
      -- 
    cr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1289_inst_req_1); -- 
    crr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => call_stmt_1203_call_req_0); -- 
    ccr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => call_stmt_1203_call_req_1); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1207_inst_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1219_inst_req_1); -- 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1229_inst_req_1); -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1239_inst_req_1); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1249_inst_req_1); -- 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1259_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1269_inst_req_1); -- 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1279_inst_req_1); -- 
    convTranspose_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(367) & convTranspose_CP_34_elements(369) & convTranspose_CP_34_elements(371) & convTranspose_CP_34_elements(373);
      gj_convTranspose_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Sample/cra
      -- 
    cra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1203_call_ack_0, ack => convTranspose_CP_34_elements(375)); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/call_stmt_1203_Update/cca
      -- CP-element group 376: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Sample/rr
      -- 
    cca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1203_call_ack_1, ack => convTranspose_CP_34_elements(376)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(376), ack => type_cast_1207_inst_req_0); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_0, ack => convTranspose_CP_34_elements(377)); -- 
    -- CP-element group 378:  fork  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	374 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	383 
    -- CP-element group 378: 	385 
    -- CP-element group 378: 	387 
    -- CP-element group 378: 	389 
    -- CP-element group 378: 	391 
    -- CP-element group 378: 	393 
    -- CP-element group 378: 	395 
    -- CP-element group 378: 	379 
    -- CP-element group 378: 	381 
    -- CP-element group 378:  members (30) 
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1207_Update/ca
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Sample/req
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Sample/rr
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_1, ack => convTranspose_CP_34_elements(378)); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1229_inst_req_0); -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1239_inst_req_0); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1249_inst_req_0); -- 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1259_inst_req_0); -- 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1269_inst_req_0); -- 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1279_inst_req_0); -- 
    rr_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1289_inst_req_0); -- 
    req_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => WPIPE_elapsed_time_pipe_1214_inst_req_0); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1219_inst_req_0); -- 
    -- CP-element group 379:  transition  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (6) 
      -- CP-element group 379: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_update_start_
      -- CP-element group 379: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Sample/ack
      -- CP-element group 379: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Update/req
      -- 
    ack_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1214_inst_ack_0, ack => convTranspose_CP_34_elements(379)); -- 
    req_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(379), ack => WPIPE_elapsed_time_pipe_1214_inst_req_1); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	420 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_elapsed_time_pipe_1214_Update/ack
      -- 
    ack_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1214_inst_ack_1, ack => convTranspose_CP_34_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	378 
    -- CP-element group 381: successors 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_0, ack => convTranspose_CP_34_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	374 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	417 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1219_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_1, ack => convTranspose_CP_34_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	378 
    -- CP-element group 383: successors 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_sample_completed_
      -- CP-element group 383: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Sample/ra
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_0, ack => convTranspose_CP_34_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	374 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	414 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_update_completed_
      -- CP-element group 384: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1229_Update/ca
      -- 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_1, ack => convTranspose_CP_34_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	378 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Sample/ra
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_0, ack => convTranspose_CP_34_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	374 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	411 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1239_Update/ca
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_1, ack => convTranspose_CP_34_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	378 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_0, ack => convTranspose_CP_34_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	374 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	408 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1249_Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_1, ack => convTranspose_CP_34_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	378 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Sample/ra
      -- 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_0, ack => convTranspose_CP_34_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	374 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	405 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1259_Update/ca
      -- 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_1, ack => convTranspose_CP_34_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	378 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Sample/ra
      -- 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_0, ack => convTranspose_CP_34_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	374 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	402 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1269_Update/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_1, ack => convTranspose_CP_34_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	378 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Sample/$exit
      -- CP-element group 393: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Sample/ra
      -- 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => convTranspose_CP_34_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	374 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	399 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Update/$exit
      -- CP-element group 394: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1279_Update/ca
      -- 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => convTranspose_CP_34_elements(394)); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	378 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Sample/ra
      -- 
    ra_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1289_inst_ack_0, ack => convTranspose_CP_34_elements(395)); -- 
    -- CP-element group 396:  transition  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	374 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (6) 
      -- CP-element group 396: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Update/ca
      -- CP-element group 396: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Sample/req
      -- CP-element group 396: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/type_cast_1289_update_completed_
      -- 
    ca_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1289_inst_ack_1, ack => convTranspose_CP_34_elements(396)); -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(396), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_0); -- 
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_update_start_
      -- CP-element group 397: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Update/req
      -- CP-element group 397: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Sample/ack
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0, ack => convTranspose_CP_34_elements(397)); -- 
    req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(397), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_1); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_update_completed_
      -- CP-element group 398: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Update/ack
      -- CP-element group 398: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1291_Update/$exit
      -- 
    ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1, ack => convTranspose_CP_34_elements(398)); -- 
    -- CP-element group 399:  join  transition  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	394 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_sample_start_
      -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(399), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_0); -- 
    convTranspose_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(394) & convTranspose_CP_34_elements(398);
      gj_convTranspose_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Update/req
      -- CP-element group 400: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Sample/ack
      -- CP-element group 400: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_update_start_
      -- CP-element group 400: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_sample_completed_
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0, ack => convTranspose_CP_34_elements(400)); -- 
    req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(400), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_1); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Update/ack
      -- CP-element group 401: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1294_update_completed_
      -- 
    ack_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1, ack => convTranspose_CP_34_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: 	392 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Sample/req
      -- CP-element group 402: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_sample_start_
      -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(402), ack => WPIPE_ConvTranspose_output_pipe_1297_inst_req_0); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(401) & convTranspose_CP_34_elements(392);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Update/req
      -- CP-element group 403: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Sample/ack
      -- CP-element group 403: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_update_start_
      -- CP-element group 403: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_sample_completed_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0, ack => convTranspose_CP_34_elements(403)); -- 
    req_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1297_inst_req_1); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Update/ack
      -- CP-element group 404: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1297_update_completed_
      -- 
    ack_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1, ack => convTranspose_CP_34_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: 	390 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Sample/req
      -- CP-element group 405: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_sample_start_
      -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(405), ack => WPIPE_ConvTranspose_output_pipe_1300_inst_req_0); -- 
    convTranspose_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(404) & convTranspose_CP_34_elements(390);
      gj_convTranspose_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Update/req
      -- CP-element group 406: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_update_start_
      -- CP-element group 406: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_sample_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0, ack => convTranspose_CP_34_elements(406)); -- 
    req_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1300_inst_req_1); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1300_update_completed_
      -- 
    ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1, ack => convTranspose_CP_34_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	388 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_sample_start_
      -- CP-element group 408: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Sample/req
      -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(408), ack => WPIPE_ConvTranspose_output_pipe_1303_inst_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(388) & convTranspose_CP_34_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Update/req
      -- CP-element group 409: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_sample_completed_
      -- CP-element group 409: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_update_start_
      -- CP-element group 409: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Sample/ack
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0, ack => convTranspose_CP_34_elements(409)); -- 
    req_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1303_inst_req_1); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1303_Update/ack
      -- 
    ack_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1, ack => convTranspose_CP_34_elements(410)); -- 
    -- CP-element group 411:  join  transition  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	386 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Sample/req
      -- CP-element group 411: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_sample_start_
      -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(411), ack => WPIPE_ConvTranspose_output_pipe_1306_inst_req_0); -- 
    convTranspose_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(386) & convTranspose_CP_34_elements(410);
      gj_convTranspose_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Update/req
      -- CP-element group 412: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_update_start_
      -- CP-element group 412: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_sample_completed_
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0, ack => convTranspose_CP_34_elements(412)); -- 
    req_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1306_inst_req_1); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1306_update_completed_
      -- 
    ack_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1, ack => convTranspose_CP_34_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	384 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_sample_start_
      -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(414), ack => WPIPE_ConvTranspose_output_pipe_1309_inst_req_0); -- 
    convTranspose_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(384) & convTranspose_CP_34_elements(413);
      gj_convTranspose_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Update/req
      -- CP-element group 415: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Sample/ack
      -- CP-element group 415: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_update_start_
      -- CP-element group 415: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_sample_completed_
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1309_inst_ack_0, ack => convTranspose_CP_34_elements(415)); -- 
    req_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1309_inst_req_1); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Update/ack
      -- CP-element group 416: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1309_update_completed_
      -- 
    ack_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1309_inst_ack_1, ack => convTranspose_CP_34_elements(416)); -- 
    -- CP-element group 417:  join  transition  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: 	382 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Sample/req
      -- CP-element group 417: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_sample_start_
      -- 
    req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(417), ack => WPIPE_ConvTranspose_output_pipe_1312_inst_req_0); -- 
    convTranspose_cp_element_group_417: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_417"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(416) & convTranspose_CP_34_elements(382);
      gj_convTranspose_cp_element_group_417 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 418:  transition  input  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (6) 
      -- CP-element group 418: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Update/req
      -- CP-element group 418: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Sample/ack
      -- CP-element group 418: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_update_start_
      -- CP-element group 418: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_sample_completed_
      -- 
    ack_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1312_inst_ack_0, ack => convTranspose_CP_34_elements(418)); -- 
    req_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(418), ack => WPIPE_ConvTranspose_output_pipe_1312_inst_req_1); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Update/ack
      -- CP-element group 419: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1312_update_completed_
      -- 
    ack_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1312_inst_ack_1, ack => convTranspose_CP_34_elements(419)); -- 
    -- CP-element group 420:  branch  join  transition  place  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: 	380 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420: 	422 
    -- CP-element group 420:  members (10) 
      -- CP-element group 420: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314__exit__
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316__entry__
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316_else_link/$entry
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316_if_link/$entry
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316_eval_test/branch_req
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316_eval_test/$exit
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316_eval_test/$entry
      -- CP-element group 420: 	 branch_block_stmt_39/if_stmt_1316_dead_link/$entry
      -- CP-element group 420: 	 branch_block_stmt_39/R_cmp264506_1317_place
      -- CP-element group 420: 	 branch_block_stmt_39/call_stmt_1203_to_assign_stmt_1314/$exit
      -- 
    branch_req_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(420), ack => if_stmt_1316_branch_req_0); -- 
    convTranspose_cp_element_group_420: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_420"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(419) & convTranspose_CP_34_elements(380);
      gj_convTranspose_cp_element_group_420 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 421:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	423 
    -- CP-element group 421: 	424 
    -- CP-element group 421:  members (18) 
      -- CP-element group 421: 	 branch_block_stmt_39/merge_stmt_1322__exit__
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357__entry__
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_update_start_
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/$entry
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_sample_start_
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Update/$entry
      -- CP-element group 421: 	 branch_block_stmt_39/if_stmt_1316_if_link/if_choice_transition
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Sample/$entry
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Sample/rr
      -- CP-element group 421: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Update/cr
      -- CP-element group 421: 	 branch_block_stmt_39/if_stmt_1316_if_link/$exit
      -- CP-element group 421: 	 branch_block_stmt_39/forx_xend273_bbx_xnph
      -- CP-element group 421: 	 branch_block_stmt_39/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 421: 	 branch_block_stmt_39/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 421: 	 branch_block_stmt_39/merge_stmt_1322_PhiReqMerge
      -- CP-element group 421: 	 branch_block_stmt_39/merge_stmt_1322_PhiAck/$entry
      -- CP-element group 421: 	 branch_block_stmt_39/merge_stmt_1322_PhiAck/$exit
      -- CP-element group 421: 	 branch_block_stmt_39/merge_stmt_1322_PhiAck/dummy
      -- 
    if_choice_transition_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1316_branch_ack_1, ack => convTranspose_CP_34_elements(421)); -- 
    rr_3112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(421), ack => type_cast_1343_inst_req_0); -- 
    cr_3117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(421), ack => type_cast_1343_inst_req_1); -- 
    -- CP-element group 422:  transition  place  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	500 
    -- CP-element group 422:  members (5) 
      -- CP-element group 422: 	 branch_block_stmt_39/if_stmt_1316_else_link/$exit
      -- CP-element group 422: 	 branch_block_stmt_39/if_stmt_1316_else_link/else_choice_transition
      -- CP-element group 422: 	 branch_block_stmt_39/forx_xend273_forx_xend501
      -- CP-element group 422: 	 branch_block_stmt_39/forx_xend273_forx_xend501_PhiReq/$entry
      -- CP-element group 422: 	 branch_block_stmt_39/forx_xend273_forx_xend501_PhiReq/$exit
      -- 
    else_choice_transition_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1316_branch_ack_0, ack => convTranspose_CP_34_elements(422)); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	421 
    -- CP-element group 423: successors 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_sample_completed_
      -- CP-element group 423: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Sample/$exit
      -- CP-element group 423: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Sample/ra
      -- 
    ra_3113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_0, ack => convTranspose_CP_34_elements(423)); -- 
    -- CP-element group 424:  transition  place  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	421 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	494 
    -- CP-element group 424:  members (9) 
      -- CP-element group 424: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357__exit__
      -- CP-element group 424: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428
      -- CP-element group 424: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/$exit
      -- CP-element group 424: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_update_completed_
      -- CP-element group 424: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Update/$exit
      -- CP-element group 424: 	 branch_block_stmt_39/assign_stmt_1328_to_assign_stmt_1357/type_cast_1343_Update/ca
      -- CP-element group 424: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/$entry
      -- CP-element group 424: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1360/$entry
      -- CP-element group 424: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/$entry
      -- 
    ca_3118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_1, ack => convTranspose_CP_34_elements(424)); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	499 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	470 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Sample/ack
      -- CP-element group 425: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_sample_complete
      -- 
    ack_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1372_index_offset_ack_0, ack => convTranspose_CP_34_elements(425)); -- 
    -- CP-element group 426:  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	499 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (11) 
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_request/req
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_request/$entry
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_base_plus_offset/sum_rename_ack
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_base_plus_offset/sum_rename_req
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_base_plus_offset/$exit
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_base_plus_offset/$entry
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Update/ack
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_offset_calculated
      -- CP-element group 426: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_root_address_calculated
      -- 
    ack_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1372_index_offset_ack_1, ack => convTranspose_CP_34_elements(426)); -- 
    req_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => addr_of_1373_final_reg_req_0); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_sample_completed_
      -- CP-element group 427: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_request/ack
      -- CP-element group 427: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_request/$exit
      -- 
    ack_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1373_final_reg_ack_0, ack => convTranspose_CP_34_elements(427)); -- 
    -- CP-element group 428:  join  fork  transition  input  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	499 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (24) 
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_plus_offset/sum_rename_ack
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_plus_offset/sum_rename_req
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_word_addrgen/$entry
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_word_addrgen/$exit
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_plus_offset/$exit
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_plus_offset/$entry
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_addr_resize/base_resize_ack
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_addr_resize/base_resize_req
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_addr_resize/$exit
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_addr_resize/$entry
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_address_resized
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_root_address_calculated
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_word_address_calculated
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_base_address_calculated
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/word_access_start/word_0/rr
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_sample_start_
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_complete/ack
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_complete/$exit
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/word_access_start/word_0/$entry
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/word_access_start/$entry
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/$entry
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_word_addrgen/root_register_ack
      -- CP-element group 428: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_word_addrgen/root_register_req
      -- 
    ack_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1373_final_reg_ack_1, ack => convTranspose_CP_34_elements(428)); -- 
    rr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(428), ack => ptr_deref_1377_load_0_req_0); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429:  members (5) 
      -- CP-element group 429: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/word_access_start/word_0/ra
      -- CP-element group 429: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/word_access_start/word_0/$exit
      -- CP-element group 429: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/word_access_start/$exit
      -- CP-element group 429: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Sample/$exit
      -- 
    ra_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1377_load_0_ack_0, ack => convTranspose_CP_34_elements(429)); -- 
    -- CP-element group 430:  fork  transition  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	499 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430: 	433 
    -- CP-element group 430: 	435 
    -- CP-element group 430: 	437 
    -- CP-element group 430: 	439 
    -- CP-element group 430: 	441 
    -- CP-element group 430: 	443 
    -- CP-element group 430: 	445 
    -- CP-element group 430:  members (33) 
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/ptr_deref_1377_Merge/merge_ack
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/ptr_deref_1377_Merge/merge_req
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/ptr_deref_1377_Merge/$exit
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/ptr_deref_1377_Merge/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/word_access_complete/word_0/ca
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/word_access_complete/word_0/$exit
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/word_access_complete/$exit
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Sample/$entry
      -- 
    ca_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1377_load_0_ack_1, ack => convTranspose_CP_34_elements(430)); -- 
    rr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1381_inst_req_0); -- 
    rr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1391_inst_req_0); -- 
    rr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1401_inst_req_0); -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1411_inst_req_0); -- 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1421_inst_req_0); -- 
    rr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1431_inst_req_0); -- 
    rr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1441_inst_req_0); -- 
    rr_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(430), ack => type_cast_1451_inst_req_0); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_sample_completed_
      -- CP-element group 431: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Sample/ra
      -- 
    ra_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_0, ack => convTranspose_CP_34_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	499 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	467 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_update_completed_
      -- CP-element group 432: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Update/ca
      -- CP-element group 432: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Update/$exit
      -- 
    ca_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_1, ack => convTranspose_CP_34_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	430 
    -- CP-element group 433: successors 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Sample/ra
      -- CP-element group 433: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Sample/$exit
      -- CP-element group 433: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_sample_completed_
      -- 
    ra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_0, ack => convTranspose_CP_34_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	499 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	464 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Update/ca
      -- CP-element group 434: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_update_completed_
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_1, ack => convTranspose_CP_34_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	430 
    -- CP-element group 435: successors 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Sample/ra
      -- CP-element group 435: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_sample_completed_
      -- 
    ra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_0, ack => convTranspose_CP_34_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	499 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	461 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_update_completed_
      -- 
    ca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_1, ack => convTranspose_CP_34_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	430 
    -- CP-element group 437: successors 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Sample/ra
      -- CP-element group 437: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Sample/$exit
      -- CP-element group 437: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_sample_completed_
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_0, ack => convTranspose_CP_34_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	499 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	458 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Update/ca
      -- CP-element group 438: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Update/$exit
      -- CP-element group 438: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_update_completed_
      -- 
    ca_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_1, ack => convTranspose_CP_34_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	430 
    -- CP-element group 439: successors 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_sample_completed_
      -- CP-element group 439: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Sample/ra
      -- CP-element group 439: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Sample/$exit
      -- 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_0, ack => convTranspose_CP_34_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	499 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	455 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_update_completed_
      -- CP-element group 440: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Update/ca
      -- CP-element group 440: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Update/$exit
      -- 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_1, ack => convTranspose_CP_34_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	430 
    -- CP-element group 441: successors 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Sample/ra
      -- CP-element group 441: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_sample_completed_
      -- 
    ra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1431_inst_ack_0, ack => convTranspose_CP_34_elements(441)); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	499 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	452 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Update/ca
      -- CP-element group 442: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_update_completed_
      -- 
    ca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1431_inst_ack_1, ack => convTranspose_CP_34_elements(442)); -- 
    -- CP-element group 443:  transition  input  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	430 
    -- CP-element group 443: successors 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Sample/ra
      -- CP-element group 443: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_sample_completed_
      -- 
    ra_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_0, ack => convTranspose_CP_34_elements(443)); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	499 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	449 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Update/ca
      -- CP-element group 444: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_update_completed_
      -- 
    ca_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_1, ack => convTranspose_CP_34_elements(444)); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	430 
    -- CP-element group 445: successors 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Sample/ra
      -- CP-element group 445: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Sample/$exit
      -- CP-element group 445: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_sample_completed_
      -- 
    ra_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1451_inst_ack_0, ack => convTranspose_CP_34_elements(445)); -- 
    -- CP-element group 446:  transition  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	499 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (6) 
      -- CP-element group 446: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Sample/req
      -- CP-element group 446: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_sample_start_
      -- CP-element group 446: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Update/ca
      -- CP-element group 446: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Update/$exit
      -- CP-element group 446: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_update_completed_
      -- 
    ca_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1451_inst_ack_1, ack => convTranspose_CP_34_elements(446)); -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1453_inst_req_0); -- 
    -- CP-element group 447:  transition  input  output  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (6) 
      -- CP-element group 447: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Update/req
      -- CP-element group 447: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Update/$entry
      -- CP-element group 447: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Sample/ack
      -- CP-element group 447: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_update_start_
      -- CP-element group 447: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_sample_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1453_inst_ack_0, ack => convTranspose_CP_34_elements(447)); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(447), ack => WPIPE_ConvTranspose_output_pipe_1453_inst_req_1); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Update/ack
      -- CP-element group 448: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1453_update_completed_
      -- 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1453_inst_ack_1, ack => convTranspose_CP_34_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	444 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Sample/req
      -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1456_inst_req_0); -- 
    convTranspose_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(444) & convTranspose_CP_34_elements(448);
      gj_convTranspose_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (6) 
      -- CP-element group 450: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Update/req
      -- CP-element group 450: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_update_start_
      -- CP-element group 450: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_sample_completed_
      -- CP-element group 450: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Sample/ack
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1456_inst_ack_0, ack => convTranspose_CP_34_elements(450)); -- 
    req_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(450), ack => WPIPE_ConvTranspose_output_pipe_1456_inst_req_1); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Update/ack
      -- CP-element group 451: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_update_completed_
      -- CP-element group 451: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1456_Update/$exit
      -- 
    ack_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1456_inst_ack_1, ack => convTranspose_CP_34_elements(451)); -- 
    -- CP-element group 452:  join  transition  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	442 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_sample_start_
      -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1459_inst_req_0); -- 
    convTranspose_cp_element_group_452: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_452"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(442) & convTranspose_CP_34_elements(451);
      gj_convTranspose_cp_element_group_452 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(452), clk => clk, reset => reset); --
    end block;
    -- CP-element group 453:  transition  input  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (6) 
      -- CP-element group 453: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Update/req
      -- CP-element group 453: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Sample/ack
      -- CP-element group 453: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Sample/$exit
      -- CP-element group 453: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_update_start_
      -- CP-element group 453: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_sample_completed_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1459_inst_ack_0, ack => convTranspose_CP_34_elements(453)); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(453), ack => WPIPE_ConvTranspose_output_pipe_1459_inst_req_1); -- 
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Update/ack
      -- CP-element group 454: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_Update/$exit
      -- CP-element group 454: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1459_update_completed_
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1459_inst_ack_1, ack => convTranspose_CP_34_elements(454)); -- 
    -- CP-element group 455:  join  transition  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	440 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_sample_start_
      -- CP-element group 455: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Sample/req
      -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1462_inst_req_0); -- 
    convTranspose_cp_element_group_455: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_455"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(440) & convTranspose_CP_34_elements(454);
      gj_convTranspose_cp_element_group_455 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 456:  transition  input  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (6) 
      -- CP-element group 456: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_sample_completed_
      -- CP-element group 456: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_update_start_
      -- CP-element group 456: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Sample/$exit
      -- CP-element group 456: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Sample/ack
      -- CP-element group 456: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Update/req
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1462_inst_ack_0, ack => convTranspose_CP_34_elements(456)); -- 
    req_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(456), ack => WPIPE_ConvTranspose_output_pipe_1462_inst_req_1); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_update_completed_
      -- CP-element group 457: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Update/$exit
      -- CP-element group 457: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1462_Update/ack
      -- 
    ack_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1462_inst_ack_1, ack => convTranspose_CP_34_elements(457)); -- 
    -- CP-element group 458:  join  transition  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	438 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_sample_start_
      -- CP-element group 458: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Sample/req
      -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1465_inst_req_0); -- 
    convTranspose_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(438) & convTranspose_CP_34_elements(457);
      gj_convTranspose_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  transition  input  output  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (6) 
      -- CP-element group 459: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_update_start_
      -- CP-element group 459: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Sample/ack
      -- CP-element group 459: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Update/$entry
      -- CP-element group 459: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Update/req
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1465_inst_ack_0, ack => convTranspose_CP_34_elements(459)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(459), ack => WPIPE_ConvTranspose_output_pipe_1465_inst_req_1); -- 
    -- CP-element group 460:  transition  input  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1465_Update/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1465_inst_ack_1, ack => convTranspose_CP_34_elements(460)); -- 
    -- CP-element group 461:  join  transition  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	436 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Sample/req
      -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1468_inst_req_0); -- 
    convTranspose_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(436) & convTranspose_CP_34_elements(460);
      gj_convTranspose_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  transition  input  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (6) 
      -- CP-element group 462: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_sample_completed_
      -- CP-element group 462: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_update_start_
      -- CP-element group 462: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Sample/$exit
      -- CP-element group 462: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Sample/ack
      -- CP-element group 462: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Update/req
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1468_inst_ack_0, ack => convTranspose_CP_34_elements(462)); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(462), ack => WPIPE_ConvTranspose_output_pipe_1468_inst_req_1); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_update_completed_
      -- CP-element group 463: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Update/$exit
      -- CP-element group 463: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1468_Update/ack
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1468_inst_ack_1, ack => convTranspose_CP_34_elements(463)); -- 
    -- CP-element group 464:  join  transition  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	434 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_sample_start_
      -- CP-element group 464: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Sample/$entry
      -- CP-element group 464: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Sample/req
      -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1471_inst_req_0); -- 
    convTranspose_cp_element_group_464: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_464"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(434) & convTranspose_CP_34_elements(463);
      gj_convTranspose_cp_element_group_464 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(464), clk => clk, reset => reset); --
    end block;
    -- CP-element group 465:  transition  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (6) 
      -- CP-element group 465: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_sample_completed_
      -- CP-element group 465: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_update_start_
      -- CP-element group 465: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Sample/$exit
      -- CP-element group 465: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Sample/ack
      -- CP-element group 465: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Update/req
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1471_inst_ack_0, ack => convTranspose_CP_34_elements(465)); -- 
    req_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(465), ack => WPIPE_ConvTranspose_output_pipe_1471_inst_req_1); -- 
    -- CP-element group 466:  transition  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Update/$exit
      -- CP-element group 466: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1471_Update/ack
      -- 
    ack_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1471_inst_ack_1, ack => convTranspose_CP_34_elements(466)); -- 
    -- CP-element group 467:  join  transition  output  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	432 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	468 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_sample_start_
      -- CP-element group 467: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Sample/$entry
      -- CP-element group 467: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Sample/req
      -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(467), ack => WPIPE_ConvTranspose_output_pipe_1474_inst_req_0); -- 
    convTranspose_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(432) & convTranspose_CP_34_elements(466);
      gj_convTranspose_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  transition  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	467 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	469 
    -- CP-element group 468:  members (6) 
      -- CP-element group 468: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_sample_completed_
      -- CP-element group 468: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_update_start_
      -- CP-element group 468: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Sample/$exit
      -- CP-element group 468: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Sample/ack
      -- CP-element group 468: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Update/req
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1474_inst_ack_0, ack => convTranspose_CP_34_elements(468)); -- 
    req_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(468), ack => WPIPE_ConvTranspose_output_pipe_1474_inst_req_1); -- 
    -- CP-element group 469:  transition  input  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	468 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	470 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_update_completed_
      -- CP-element group 469: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Update/$exit
      -- CP-element group 469: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/WPIPE_ConvTranspose_output_pipe_1474_Update/ack
      -- 
    ack_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1474_inst_ack_1, ack => convTranspose_CP_34_elements(469)); -- 
    -- CP-element group 470:  branch  join  transition  place  output  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	425 
    -- CP-element group 470: 	469 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470: 	472 
    -- CP-element group 470:  members (10) 
      -- CP-element group 470: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487__exit__
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488__entry__
      -- CP-element group 470: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/$exit
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488_dead_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488_eval_test/$entry
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488_eval_test/$exit
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488_eval_test/branch_req
      -- CP-element group 470: 	 branch_block_stmt_39/R_exitcond1_1489_place
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488_if_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_39/if_stmt_1488_else_link/$entry
      -- 
    branch_req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(470), ack => if_stmt_1488_branch_req_0); -- 
    convTranspose_cp_element_group_470: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_470"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(425) & convTranspose_CP_34_elements(469);
      gj_convTranspose_cp_element_group_470 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(470), clk => clk, reset => reset); --
    end block;
    -- CP-element group 471:  merge  transition  place  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	470 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	500 
    -- CP-element group 471:  members (13) 
      -- CP-element group 471: 	 branch_block_stmt_39/merge_stmt_1494__exit__
      -- CP-element group 471: 	 branch_block_stmt_39/forx_xend501x_xloopexit_forx_xend501
      -- CP-element group 471: 	 branch_block_stmt_39/if_stmt_1488_if_link/$exit
      -- CP-element group 471: 	 branch_block_stmt_39/if_stmt_1488_if_link/if_choice_transition
      -- CP-element group 471: 	 branch_block_stmt_39/forx_xbody428_forx_xend501x_xloopexit
      -- CP-element group 471: 	 branch_block_stmt_39/forx_xbody428_forx_xend501x_xloopexit_PhiReq/$entry
      -- CP-element group 471: 	 branch_block_stmt_39/forx_xbody428_forx_xend501x_xloopexit_PhiReq/$exit
      -- CP-element group 471: 	 branch_block_stmt_39/merge_stmt_1494_PhiReqMerge
      -- CP-element group 471: 	 branch_block_stmt_39/merge_stmt_1494_PhiAck/$entry
      -- CP-element group 471: 	 branch_block_stmt_39/merge_stmt_1494_PhiAck/$exit
      -- CP-element group 471: 	 branch_block_stmt_39/merge_stmt_1494_PhiAck/dummy
      -- CP-element group 471: 	 branch_block_stmt_39/forx_xend501x_xloopexit_forx_xend501_PhiReq/$entry
      -- CP-element group 471: 	 branch_block_stmt_39/forx_xend501x_xloopexit_forx_xend501_PhiReq/$exit
      -- 
    if_choice_transition_3454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_1, ack => convTranspose_CP_34_elements(471)); -- 
    -- CP-element group 472:  fork  transition  place  input  output  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	470 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	495 
    -- CP-element group 472: 	496 
    -- CP-element group 472:  members (12) 
      -- CP-element group 472: 	 branch_block_stmt_39/if_stmt_1488_else_link/$exit
      -- CP-element group 472: 	 branch_block_stmt_39/if_stmt_1488_else_link/else_choice_transition
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Sample/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Sample/rr
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Update/$entry
      -- CP-element group 472: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_0, ack => convTranspose_CP_34_elements(472)); -- 
    rr_3733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(472), ack => type_cast_1366_inst_req_0); -- 
    cr_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(472), ack => type_cast_1366_inst_req_1); -- 
    -- CP-element group 473:  merge  branch  transition  place  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	165 
    -- CP-element group 473: 	120 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	121 
    -- CP-element group 473: 	122 
    -- CP-element group 473:  members (17) 
      -- CP-element group 473: 	 branch_block_stmt_39/merge_stmt_430__exit__
      -- CP-element group 473: 	 branch_block_stmt_39/assign_stmt_436__entry__
      -- CP-element group 473: 	 branch_block_stmt_39/assign_stmt_436__exit__
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437__entry__
      -- CP-element group 473: 	 branch_block_stmt_39/assign_stmt_436/$entry
      -- CP-element group 473: 	 branch_block_stmt_39/assign_stmt_436/$exit
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437_dead_link/$entry
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437_eval_test/$entry
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437_eval_test/$exit
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437_eval_test/branch_req
      -- CP-element group 473: 	 branch_block_stmt_39/R_cmp194510_438_place
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437_if_link/$entry
      -- CP-element group 473: 	 branch_block_stmt_39/if_stmt_437_else_link/$entry
      -- CP-element group 473: 	 branch_block_stmt_39/merge_stmt_430_PhiReqMerge
      -- CP-element group 473: 	 branch_block_stmt_39/merge_stmt_430_PhiAck/$entry
      -- CP-element group 473: 	 branch_block_stmt_39/merge_stmt_430_PhiAck/$exit
      -- CP-element group 473: 	 branch_block_stmt_39/merge_stmt_430_PhiAck/dummy
      -- 
    branch_req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(473), ack => if_stmt_437_branch_req_0); -- 
    convTranspose_CP_34_elements(473) <= OrReduce(convTranspose_CP_34_elements(165) & convTranspose_CP_34_elements(120));
    -- CP-element group 474:  transition  output  delay-element  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	124 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	478 
    -- CP-element group 474:  members (5) 
      -- CP-element group 474: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/$exit
      -- CP-element group 474: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_475/$exit
      -- CP-element group 474: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/$exit
      -- CP-element group 474: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_479_konst_delay_trans
      -- CP-element group 474: 	 branch_block_stmt_39/bbx_xnph516_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_req
      -- 
    phi_stmt_475_req_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_475_req_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(474), ack => phi_stmt_475_req_0); -- 
    -- Element group convTranspose_CP_34_elements(474) is a control-delay.
    cp_element_474_delay: control_delay_element  generic map(name => " 474_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(124), ack => convTranspose_CP_34_elements(474), clk => clk, reset =>reset);
    -- CP-element group 475:  transition  input  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	166 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	477 
    -- CP-element group 475:  members (2) 
      -- CP-element group 475: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Sample/$exit
      -- CP-element group 475: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Sample/ra
      -- 
    ra_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_0, ack => convTranspose_CP_34_elements(475)); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	166 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	477 
    -- CP-element group 476:  members (2) 
      -- CP-element group 476: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Update/$exit
      -- CP-element group 476: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/Update/ca
      -- 
    ca_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_1, ack => convTranspose_CP_34_elements(476)); -- 
    -- CP-element group 477:  join  transition  output  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	475 
    -- CP-element group 477: 	476 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	478 
    -- CP-element group 477:  members (6) 
      -- CP-element group 477: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 477: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/$exit
      -- CP-element group 477: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/$exit
      -- CP-element group 477: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/$exit
      -- CP-element group 477: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_sources/type_cast_481/SplitProtocol/$exit
      -- CP-element group 477: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_475/phi_stmt_475_req
      -- 
    phi_stmt_475_req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_475_req_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(477), ack => phi_stmt_475_req_1); -- 
    convTranspose_cp_element_group_477: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_477"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(475) & convTranspose_CP_34_elements(476);
      gj_convTranspose_cp_element_group_477 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 478:  merge  transition  place  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	474 
    -- CP-element group 478: 	477 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	479 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_39/merge_stmt_474_PhiReqMerge
      -- CP-element group 478: 	 branch_block_stmt_39/merge_stmt_474_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(478) <= OrReduce(convTranspose_CP_34_elements(474) & convTranspose_CP_34_elements(477));
    -- CP-element group 479:  fork  transition  place  input  output  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	478 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	163 
    -- CP-element group 479: 	125 
    -- CP-element group 479: 	126 
    -- CP-element group 479: 	128 
    -- CP-element group 479: 	129 
    -- CP-element group 479: 	132 
    -- CP-element group 479: 	136 
    -- CP-element group 479: 	140 
    -- CP-element group 479: 	144 
    -- CP-element group 479: 	148 
    -- CP-element group 479: 	152 
    -- CP-element group 479: 	156 
    -- CP-element group 479: 	160 
    -- CP-element group 479:  members (56) 
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/merge_stmt_474__exit__
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637__entry__
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_544_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_598_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/word_access_complete/word_0/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/word_access_complete/word_0/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/word_access_complete/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_580_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_616_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_562_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/ptr_deref_624_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_resized_1
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_scaled_1
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_computed_1
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_resize_1/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_resize_1/$exit
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_resize_1/index_resize_req
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_resize_1/index_resize_ack
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_scale_1/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_scale_1/$exit
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_scale_1/scale_rename_req
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_index_scale_1/scale_rename_ack
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_update_start
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Sample/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Sample/req
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/array_obj_ref_487_final_index_sum_regn_Update/req
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_complete/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/addr_of_488_complete/req
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_sample_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Sample/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/RPIPE_ConvTranspose_input_pipe_491_Sample/rr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_495_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_508_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_update_start_
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_39/assign_stmt_489_to_assign_stmt_637/type_cast_526_Update/cr
      -- CP-element group 479: 	 branch_block_stmt_39/merge_stmt_474_PhiAck/$exit
      -- CP-element group 479: 	 branch_block_stmt_39/merge_stmt_474_PhiAck/phi_stmt_475_ack
      -- 
    phi_stmt_475_ack_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_475_ack_0, ack => convTranspose_CP_34_elements(479)); -- 
    cr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_544_inst_req_1); -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_598_inst_req_1); -- 
    cr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => ptr_deref_624_store_0_req_1); -- 
    cr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_616_inst_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_580_inst_req_1); -- 
    cr_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_562_inst_req_1); -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => array_obj_ref_487_index_offset_req_0); -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => array_obj_ref_487_index_offset_req_1); -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => addr_of_488_final_reg_req_1); -- 
    rr_1009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => RPIPE_ConvTranspose_input_pipe_491_inst_req_0); -- 
    cr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_495_inst_req_1); -- 
    cr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_508_inst_req_1); -- 
    cr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => type_cast_526_inst_req_1); -- 
    -- CP-element group 480:  transition  output  delay-element  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	168 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	484 
    -- CP-element group 480:  members (5) 
      -- CP-element group 480: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/$exit
      -- CP-element group 480: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_682/$exit
      -- CP-element group 480: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/$exit
      -- CP-element group 480: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_688_konst_delay_trans
      -- CP-element group 480: 	 branch_block_stmt_39/bbx_xnph512_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_req
      -- 
    phi_stmt_682_req_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_682_req_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(480), ack => phi_stmt_682_req_1); -- 
    -- Element group convTranspose_CP_34_elements(480) is a control-delay.
    cp_element_480_delay: control_delay_element  generic map(name => " 480_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(168), ack => convTranspose_CP_34_elements(480), clk => clk, reset =>reset);
    -- CP-element group 481:  transition  input  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	210 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	483 
    -- CP-element group 481:  members (2) 
      -- CP-element group 481: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Sample/$exit
      -- CP-element group 481: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Sample/ra
      -- 
    ra_3580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_685_inst_ack_0, ack => convTranspose_CP_34_elements(481)); -- 
    -- CP-element group 482:  transition  input  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	210 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482:  members (2) 
      -- CP-element group 482: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Update/$exit
      -- CP-element group 482: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/Update/ca
      -- 
    ca_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_685_inst_ack_1, ack => convTranspose_CP_34_elements(482)); -- 
    -- CP-element group 483:  join  transition  output  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	481 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	484 
    -- CP-element group 483:  members (6) 
      -- CP-element group 483: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 483: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/$exit
      -- CP-element group 483: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/$exit
      -- CP-element group 483: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/$exit
      -- CP-element group 483: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_sources/type_cast_685/SplitProtocol/$exit
      -- CP-element group 483: 	 branch_block_stmt_39/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_682/phi_stmt_682_req
      -- 
    phi_stmt_682_req_3586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_682_req_3586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => phi_stmt_682_req_0); -- 
    convTranspose_cp_element_group_483: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_483"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(481) & convTranspose_CP_34_elements(482);
      gj_convTranspose_cp_element_group_483 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(483), clk => clk, reset => reset); --
    end block;
    -- CP-element group 484:  merge  transition  place  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	480 
    -- CP-element group 484: 	483 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	485 
    -- CP-element group 484:  members (2) 
      -- CP-element group 484: 	 branch_block_stmt_39/merge_stmt_681_PhiReqMerge
      -- CP-element group 484: 	 branch_block_stmt_39/merge_stmt_681_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(484) <= OrReduce(convTranspose_CP_34_elements(480) & convTranspose_CP_34_elements(483));
    -- CP-element group 485:  fork  transition  place  input  output  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	484 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	184 
    -- CP-element group 485: 	188 
    -- CP-element group 485: 	192 
    -- CP-element group 485: 	196 
    -- CP-element group 485: 	200 
    -- CP-element group 485: 	204 
    -- CP-element group 485: 	207 
    -- CP-element group 485: 	180 
    -- CP-element group 485: 	169 
    -- CP-element group 485: 	170 
    -- CP-element group 485: 	172 
    -- CP-element group 485: 	173 
    -- CP-element group 485: 	176 
    -- CP-element group 485:  members (56) 
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_complete/req
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_complete/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/merge_stmt_681__exit__
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844__entry__
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/addr_of_695_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_sample_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Update/req
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Sample/req
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_733_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Sample/rr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_final_index_sum_regn_update_start
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_715_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/RPIPE_ConvTranspose_input_pipe_698_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_scale_1/scale_rename_ack
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_702_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_scale_1/scale_rename_req
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_scale_1/$exit
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_scale_1/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_resize_1/index_resize_ack
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_resize_1/index_resize_req
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_resize_1/$exit
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_resize_1/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_computed_1
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_scaled_1
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/array_obj_ref_694_index_resized_1
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_751_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_769_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_787_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_805_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/type_cast_823_Update/cr
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_update_start_
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/word_access_complete/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/word_access_complete/word_0/$entry
      -- CP-element group 485: 	 branch_block_stmt_39/assign_stmt_696_to_assign_stmt_844/ptr_deref_831_Update/word_access_complete/word_0/cr
      -- CP-element group 485: 	 branch_block_stmt_39/merge_stmt_681_PhiAck/$exit
      -- CP-element group 485: 	 branch_block_stmt_39/merge_stmt_681_PhiAck/phi_stmt_682_ack
      -- 
    phi_stmt_682_ack_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_682_ack_0, ack => convTranspose_CP_34_elements(485)); -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => addr_of_695_final_reg_req_1); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => array_obj_ref_694_index_offset_req_1); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => array_obj_ref_694_index_offset_req_0); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_715_inst_req_1); -- 
    cr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_733_inst_req_1); -- 
    rr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => RPIPE_ConvTranspose_input_pipe_698_inst_req_0); -- 
    cr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_702_inst_req_1); -- 
    cr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_751_inst_req_1); -- 
    cr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_769_inst_req_1); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_787_inst_req_1); -- 
    cr_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_805_inst_req_1); -- 
    cr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => type_cast_823_inst_req_1); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(485), ack => ptr_deref_831_store_0_req_1); -- 
    -- CP-element group 486:  merge  fork  transition  place  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	209 
    -- CP-element group 486: 	122 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	211 
    -- CP-element group 486: 	212 
    -- CP-element group 486: 	213 
    -- CP-element group 486: 	214 
    -- CP-element group 486: 	215 
    -- CP-element group 486: 	216 
    -- CP-element group 486:  members (25) 
      -- CP-element group 486: 	 branch_block_stmt_39/merge_stmt_853__exit__
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881__entry__
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_update_start_
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Sample/rr
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Update/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_856_Update/cr
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_update_start_
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Sample/rr
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Update/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_860_Update/cr
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_update_start_
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Sample/rr
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Update/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/assign_stmt_857_to_assign_stmt_881/type_cast_864_Update/cr
      -- CP-element group 486: 	 branch_block_stmt_39/merge_stmt_853_PhiReqMerge
      -- CP-element group 486: 	 branch_block_stmt_39/merge_stmt_853_PhiAck/$entry
      -- CP-element group 486: 	 branch_block_stmt_39/merge_stmt_853_PhiAck/$exit
      -- CP-element group 486: 	 branch_block_stmt_39/merge_stmt_853_PhiAck/dummy
      -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => type_cast_856_inst_req_0); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => type_cast_856_inst_req_1); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => type_cast_860_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => type_cast_860_inst_req_1); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => type_cast_864_inst_req_0); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => type_cast_864_inst_req_1); -- 
    convTranspose_CP_34_elements(486) <= OrReduce(convTranspose_CP_34_elements(209) & convTranspose_CP_34_elements(122));
    -- CP-element group 487:  transition  output  delay-element  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	221 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	491 
    -- CP-element group 487:  members (5) 
      -- CP-element group 487: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/$exit
      -- CP-element group 487: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_926/$exit
      -- CP-element group 487: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/$exit
      -- CP-element group 487: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_932_konst_delay_trans
      -- CP-element group 487: 	 branch_block_stmt_39/bbx_xnph508_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_req
      -- 
    phi_stmt_926_req_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_926_req_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(487), ack => phi_stmt_926_req_1); -- 
    -- Element group convTranspose_CP_34_elements(487) is a control-delay.
    cp_element_487_delay: control_delay_element  generic map(name => " 487_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(221), ack => convTranspose_CP_34_elements(487), clk => clk, reset =>reset);
    -- CP-element group 488:  transition  input  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	230 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	490 
    -- CP-element group 488:  members (2) 
      -- CP-element group 488: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Sample/$exit
      -- CP-element group 488: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Sample/ra
      -- 
    ra_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_929_inst_ack_0, ack => convTranspose_CP_34_elements(488)); -- 
    -- CP-element group 489:  transition  input  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	230 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489:  members (2) 
      -- CP-element group 489: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Update/$exit
      -- CP-element group 489: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/Update/ca
      -- 
    ca_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_929_inst_ack_1, ack => convTranspose_CP_34_elements(489)); -- 
    -- CP-element group 490:  join  transition  output  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	488 
    -- CP-element group 490: 	489 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (6) 
      -- CP-element group 490: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 490: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/$exit
      -- CP-element group 490: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/$exit
      -- CP-element group 490: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/$exit
      -- CP-element group 490: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_sources/type_cast_929/SplitProtocol/$exit
      -- CP-element group 490: 	 branch_block_stmt_39/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_926/phi_stmt_926_req
      -- 
    phi_stmt_926_req_3663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_926_req_3663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => phi_stmt_926_req_0); -- 
    convTranspose_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(488) & convTranspose_CP_34_elements(489);
      gj_convTranspose_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  merge  transition  place  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	487 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	492 
    -- CP-element group 491:  members (2) 
      -- CP-element group 491: 	 branch_block_stmt_39/merge_stmt_925_PhiReqMerge
      -- CP-element group 491: 	 branch_block_stmt_39/merge_stmt_925_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(491) <= OrReduce(convTranspose_CP_34_elements(487) & convTranspose_CP_34_elements(490));
    -- CP-element group 492:  fork  transition  place  input  output  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	491 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	222 
    -- CP-element group 492: 	223 
    -- CP-element group 492: 	225 
    -- CP-element group 492: 	227 
    -- CP-element group 492:  members (29) 
      -- CP-element group 492: 	 branch_block_stmt_39/merge_stmt_925__exit__
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956__entry__
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_update_start_
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_resized_1
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_scaled_1
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_computed_1
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_resize_1/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_resize_1/$exit
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_resize_1/index_resize_req
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_resize_1/index_resize_ack
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_scale_1/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_scale_1/$exit
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_scale_1/scale_rename_req
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_index_scale_1/scale_rename_ack
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_update_start
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Sample/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Sample/req
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Update/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/array_obj_ref_938_final_index_sum_regn_Update/req
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_complete/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/addr_of_939_complete/req
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_update_start_
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/word_access_complete/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/word_access_complete/word_0/$entry
      -- CP-element group 492: 	 branch_block_stmt_39/assign_stmt_940_to_assign_stmt_956/ptr_deref_942_Update/word_access_complete/word_0/cr
      -- CP-element group 492: 	 branch_block_stmt_39/merge_stmt_925_PhiAck/$exit
      -- CP-element group 492: 	 branch_block_stmt_39/merge_stmt_925_PhiAck/phi_stmt_926_ack
      -- 
    phi_stmt_926_ack_3668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_926_ack_0, ack => convTranspose_CP_34_elements(492)); -- 
    req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(492), ack => array_obj_ref_938_index_offset_req_0); -- 
    req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(492), ack => array_obj_ref_938_index_offset_req_1); -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(492), ack => addr_of_939_final_reg_req_1); -- 
    cr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(492), ack => ptr_deref_942_store_0_req_1); -- 
    -- CP-element group 493:  merge  fork  transition  place  output  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	219 
    -- CP-element group 493: 	229 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	231 
    -- CP-element group 493: 	232 
    -- CP-element group 493: 	234 
    -- CP-element group 493:  members (16) 
      -- CP-element group 493: 	 branch_block_stmt_39/merge_stmt_965__exit__
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974__entry__
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/$entry
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_sample_start_
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_update_start_
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Sample/$entry
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Sample/crr
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Update/$entry
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/call_stmt_968_Update/ccr
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_update_start_
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Update/$entry
      -- CP-element group 493: 	 branch_block_stmt_39/call_stmt_968_to_assign_stmt_974/type_cast_973_Update/cr
      -- CP-element group 493: 	 branch_block_stmt_39/merge_stmt_965_PhiReqMerge
      -- CP-element group 493: 	 branch_block_stmt_39/merge_stmt_965_PhiAck/$entry
      -- CP-element group 493: 	 branch_block_stmt_39/merge_stmt_965_PhiAck/$exit
      -- CP-element group 493: 	 branch_block_stmt_39/merge_stmt_965_PhiAck/dummy
      -- 
    crr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(493), ack => call_stmt_968_call_req_0); -- 
    ccr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(493), ack => call_stmt_968_call_req_1); -- 
    cr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(493), ack => type_cast_973_inst_req_1); -- 
    convTranspose_CP_34_elements(493) <= OrReduce(convTranspose_CP_34_elements(219) & convTranspose_CP_34_elements(229));
    -- CP-element group 494:  transition  output  delay-element  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	424 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	498 
    -- CP-element group 494:  members (5) 
      -- CP-element group 494: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/$exit
      -- CP-element group 494: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1360/$exit
      -- CP-element group 494: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/$exit
      -- CP-element group 494: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1364_konst_delay_trans
      -- CP-element group 494: 	 branch_block_stmt_39/bbx_xnph_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_req
      -- 
    phi_stmt_1360_req_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1360_req_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(494), ack => phi_stmt_1360_req_0); -- 
    -- Element group convTranspose_CP_34_elements(494) is a control-delay.
    cp_element_494_delay: control_delay_element  generic map(name => " 494_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(424), ack => convTranspose_CP_34_elements(494), clk => clk, reset =>reset);
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	472 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	497 
    -- CP-element group 495:  members (2) 
      -- CP-element group 495: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Sample/$exit
      -- CP-element group 495: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Sample/ra
      -- 
    ra_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => convTranspose_CP_34_elements(495)); -- 
    -- CP-element group 496:  transition  input  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	472 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (2) 
      -- CP-element group 496: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Update/$exit
      -- CP-element group 496: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/Update/ca
      -- 
    ca_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => convTranspose_CP_34_elements(496)); -- 
    -- CP-element group 497:  join  transition  output  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	495 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (6) 
      -- CP-element group 497: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/$exit
      -- CP-element group 497: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/$exit
      -- CP-element group 497: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/$exit
      -- CP-element group 497: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/$exit
      -- CP-element group 497: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_sources/type_cast_1366/SplitProtocol/$exit
      -- CP-element group 497: 	 branch_block_stmt_39/forx_xbody428_forx_xbody428_PhiReq/phi_stmt_1360/phi_stmt_1360_req
      -- 
    phi_stmt_1360_req_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1360_req_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(497), ack => phi_stmt_1360_req_1); -- 
    convTranspose_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(495) & convTranspose_CP_34_elements(496);
      gj_convTranspose_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  merge  transition  place  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	494 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	499 
    -- CP-element group 498:  members (2) 
      -- CP-element group 498: 	 branch_block_stmt_39/merge_stmt_1359_PhiReqMerge
      -- CP-element group 498: 	 branch_block_stmt_39/merge_stmt_1359_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(498) <= OrReduce(convTranspose_CP_34_elements(494) & convTranspose_CP_34_elements(497));
    -- CP-element group 499:  fork  transition  place  input  output  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	498 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	425 
    -- CP-element group 499: 	426 
    -- CP-element group 499: 	428 
    -- CP-element group 499: 	430 
    -- CP-element group 499: 	432 
    -- CP-element group 499: 	434 
    -- CP-element group 499: 	436 
    -- CP-element group 499: 	438 
    -- CP-element group 499: 	440 
    -- CP-element group 499: 	442 
    -- CP-element group 499: 	444 
    -- CP-element group 499: 	446 
    -- CP-element group 499:  members (53) 
      -- CP-element group 499: 	 branch_block_stmt_39/merge_stmt_1359__exit__
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487__entry__
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1401_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/word_access_complete/word_0/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/word_access_complete/word_0/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/word_access_complete/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/ptr_deref_1377_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_complete/req
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/addr_of_1373_complete/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1451_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Update/req
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1391_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Sample/req
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1441_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_final_index_sum_regn_update_start
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_scale_1/scale_rename_ack
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_scale_1/scale_rename_req
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_scale_1/$exit
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_scale_1/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_resize_1/index_resize_ack
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1411_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_resize_1/index_resize_req
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_resize_1/$exit
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_resize_1/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1431_update_start_
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_computed_1
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Update/cr
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1381_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_scaled_1
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/array_obj_ref_1372_index_resized_1
      -- CP-element group 499: 	 branch_block_stmt_39/assign_stmt_1374_to_assign_stmt_1487/type_cast_1421_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_39/merge_stmt_1359_PhiAck/$exit
      -- CP-element group 499: 	 branch_block_stmt_39/merge_stmt_1359_PhiAck/phi_stmt_1360_ack
      -- 
    phi_stmt_1360_ack_3745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1360_ack_0, ack => convTranspose_CP_34_elements(499)); -- 
    cr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1401_inst_req_1); -- 
    cr_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1411_inst_req_1); -- 
    cr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => ptr_deref_1377_load_0_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1391_inst_req_1); -- 
    req_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => addr_of_1373_final_reg_req_1); -- 
    cr_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1451_inst_req_1); -- 
    req_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => array_obj_ref_1372_index_offset_req_1); -- 
    cr_3314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1441_inst_req_1); -- 
    req_3146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => array_obj_ref_1372_index_offset_req_0); -- 
    cr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1431_inst_req_1); -- 
    cr_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1381_inst_req_1); -- 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(499), ack => type_cast_1421_inst_req_1); -- 
    -- CP-element group 500:  merge  transition  place  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	422 
    -- CP-element group 500: 	471 
    -- CP-element group 500: successors 
    -- CP-element group 500:  members (16) 
      -- CP-element group 500: 	 $exit
      -- CP-element group 500: 	 branch_block_stmt_39/$exit
      -- CP-element group 500: 	 branch_block_stmt_39/branch_block_stmt_39__exit__
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1496__exit__
      -- CP-element group 500: 	 branch_block_stmt_39/return__
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1498__exit__
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1496_PhiReqMerge
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1496_PhiAck/$entry
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1496_PhiAck/$exit
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1496_PhiAck/dummy
      -- CP-element group 500: 	 branch_block_stmt_39/return___PhiReq/$entry
      -- CP-element group 500: 	 branch_block_stmt_39/return___PhiReq/$exit
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1498_PhiReqMerge
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1498_PhiAck/$entry
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1498_PhiAck/$exit
      -- CP-element group 500: 	 branch_block_stmt_39/merge_stmt_1498_PhiAck/dummy
      -- 
    convTranspose_CP_34_elements(500) <= OrReduce(convTranspose_CP_34_elements(422) & convTranspose_CP_34_elements(471));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar526_937_resized : std_logic_vector(13 downto 0);
    signal R_indvar526_937_scaled : std_logic_vector(13 downto 0);
    signal R_indvar540_693_resized : std_logic_vector(10 downto 0);
    signal R_indvar540_693_scaled : std_logic_vector(10 downto 0);
    signal R_indvar556_486_resized : std_logic_vector(13 downto 0);
    signal R_indvar556_486_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1371_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1371_scaled : std_logic_vector(13 downto 0);
    signal add108_340 : std_logic_vector(15 downto 0);
    signal add117_365 : std_logic_vector(15 downto 0);
    signal add126_390 : std_logic_vector(15 downto 0);
    signal add12_89 : std_logic_vector(15 downto 0);
    signal add135_415 : std_logic_vector(15 downto 0);
    signal add150_514 : std_logic_vector(63 downto 0);
    signal add156_532 : std_logic_vector(63 downto 0);
    signal add162_550 : std_logic_vector(63 downto 0);
    signal add168_568 : std_logic_vector(63 downto 0);
    signal add174_586 : std_logic_vector(63 downto 0);
    signal add180_604 : std_logic_vector(63 downto 0);
    signal add186_622 : std_logic_vector(63 downto 0);
    signal add206_721 : std_logic_vector(63 downto 0);
    signal add212_739 : std_logic_vector(63 downto 0);
    signal add218_757 : std_logic_vector(63 downto 0);
    signal add21_114 : std_logic_vector(15 downto 0);
    signal add224_775 : std_logic_vector(63 downto 0);
    signal add230_793 : std_logic_vector(63 downto 0);
    signal add236_811 : std_logic_vector(63 downto 0);
    signal add242_829 : std_logic_vector(63 downto 0);
    signal add30_139 : std_logic_vector(15 downto 0);
    signal add39_164 : std_logic_vector(15 downto 0);
    signal add48_189 : std_logic_vector(15 downto 0);
    signal add57_214 : std_logic_vector(15 downto 0);
    signal add74_254 : std_logic_vector(31 downto 0);
    signal add79_259 : std_logic_vector(31 downto 0);
    signal add99_315 : std_logic_vector(15 downto 0);
    signal add_64 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1372_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1372_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1372_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1372_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1372_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1372_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_487_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_487_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_487_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_487_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_487_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_487_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_694_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_694_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_694_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_694_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_694_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_694_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_938_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_938_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_938_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_938_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_938_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_938_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_696 : std_logic_vector(31 downto 0);
    signal arrayidx269_940 : std_logic_vector(31 downto 0);
    signal arrayidx433_1374 : std_logic_vector(31 downto 0);
    signal arrayidx_489 : std_logic_vector(31 downto 0);
    signal call101_318 : std_logic_vector(7 downto 0);
    signal call106_331 : std_logic_vector(7 downto 0);
    signal call10_80 : std_logic_vector(7 downto 0);
    signal call110_343 : std_logic_vector(7 downto 0);
    signal call115_356 : std_logic_vector(7 downto 0);
    signal call119_368 : std_logic_vector(7 downto 0);
    signal call124_381 : std_logic_vector(7 downto 0);
    signal call128_393 : std_logic_vector(7 downto 0);
    signal call133_406 : std_logic_vector(7 downto 0);
    signal call143_492 : std_logic_vector(7 downto 0);
    signal call147_505 : std_logic_vector(7 downto 0);
    signal call14_92 : std_logic_vector(7 downto 0);
    signal call153_523 : std_logic_vector(7 downto 0);
    signal call159_541 : std_logic_vector(7 downto 0);
    signal call165_559 : std_logic_vector(7 downto 0);
    signal call171_577 : std_logic_vector(7 downto 0);
    signal call177_595 : std_logic_vector(7 downto 0);
    signal call183_613 : std_logic_vector(7 downto 0);
    signal call199_699 : std_logic_vector(7 downto 0);
    signal call19_105 : std_logic_vector(7 downto 0);
    signal call203_712 : std_logic_vector(7 downto 0);
    signal call209_730 : std_logic_vector(7 downto 0);
    signal call215_748 : std_logic_vector(7 downto 0);
    signal call221_766 : std_logic_vector(7 downto 0);
    signal call227_784 : std_logic_vector(7 downto 0);
    signal call233_802 : std_logic_vector(7 downto 0);
    signal call239_820 : std_logic_vector(7 downto 0);
    signal call23_117 : std_logic_vector(7 downto 0);
    signal call275_968 : std_logic_vector(63 downto 0);
    signal call28_130 : std_logic_vector(7 downto 0);
    signal call2_55 : std_logic_vector(7 downto 0);
    signal call32_142 : std_logic_vector(7 downto 0);
    signal call346_1191 : std_logic_vector(15 downto 0);
    signal call348_1194 : std_logic_vector(15 downto 0);
    signal call350_1197 : std_logic_vector(15 downto 0);
    signal call352_1200 : std_logic_vector(15 downto 0);
    signal call354_1203 : std_logic_vector(63 downto 0);
    signal call37_155 : std_logic_vector(7 downto 0);
    signal call41_167 : std_logic_vector(7 downto 0);
    signal call46_180 : std_logic_vector(7 downto 0);
    signal call50_192 : std_logic_vector(7 downto 0);
    signal call55_205 : std_logic_vector(7 downto 0);
    signal call5_67 : std_logic_vector(7 downto 0);
    signal call92_293 : std_logic_vector(7 downto 0);
    signal call97_306 : std_logic_vector(7 downto 0);
    signal call_42 : std_logic_vector(7 downto 0);
    signal cmp194510_436 : std_logic_vector(0 downto 0);
    signal cmp264506_881 : std_logic_vector(0 downto 0);
    signal cmp514_421 : std_logic_vector(0 downto 0);
    signal conv104_322 : std_logic_vector(15 downto 0);
    signal conv107_335 : std_logic_vector(15 downto 0);
    signal conv113_347 : std_logic_vector(15 downto 0);
    signal conv116_360 : std_logic_vector(15 downto 0);
    signal conv11_84 : std_logic_vector(15 downto 0);
    signal conv122_372 : std_logic_vector(15 downto 0);
    signal conv125_385 : std_logic_vector(15 downto 0);
    signal conv131_397 : std_logic_vector(15 downto 0);
    signal conv134_410 : std_logic_vector(15 downto 0);
    signal conv144_496 : std_logic_vector(63 downto 0);
    signal conv149_509 : std_logic_vector(63 downto 0);
    signal conv155_527 : std_logic_vector(63 downto 0);
    signal conv161_545 : std_logic_vector(63 downto 0);
    signal conv167_563 : std_logic_vector(63 downto 0);
    signal conv173_581 : std_logic_vector(63 downto 0);
    signal conv179_599 : std_logic_vector(63 downto 0);
    signal conv17_96 : std_logic_vector(15 downto 0);
    signal conv185_617 : std_logic_vector(63 downto 0);
    signal conv1_46 : std_logic_vector(15 downto 0);
    signal conv200_703 : std_logic_vector(63 downto 0);
    signal conv205_716 : std_logic_vector(63 downto 0);
    signal conv20_109 : std_logic_vector(15 downto 0);
    signal conv211_734 : std_logic_vector(63 downto 0);
    signal conv217_752 : std_logic_vector(63 downto 0);
    signal conv223_770 : std_logic_vector(63 downto 0);
    signal conv229_788 : std_logic_vector(63 downto 0);
    signal conv235_806 : std_logic_vector(63 downto 0);
    signal conv241_824 : std_logic_vector(63 downto 0);
    signal conv253_857 : std_logic_vector(31 downto 0);
    signal conv255_861 : std_logic_vector(31 downto 0);
    signal conv258_865 : std_logic_vector(31 downto 0);
    signal conv26_121 : std_logic_vector(15 downto 0);
    signal conv276_974 : std_logic_vector(63 downto 0);
    signal conv29_134 : std_logic_vector(15 downto 0);
    signal conv305_1056 : std_logic_vector(15 downto 0);
    signal conv307_1063 : std_logic_vector(15 downto 0);
    signal conv322_1112 : std_logic_vector(15 downto 0);
    signal conv324_1119 : std_logic_vector(15 downto 0);
    signal conv339_1168 : std_logic_vector(15 downto 0);
    signal conv341_1175 : std_logic_vector(15 downto 0);
    signal conv355_1208 : std_logic_vector(63 downto 0);
    signal conv35_146 : std_logic_vector(15 downto 0);
    signal conv362_1220 : std_logic_vector(7 downto 0);
    signal conv368_1230 : std_logic_vector(7 downto 0);
    signal conv374_1240 : std_logic_vector(7 downto 0);
    signal conv380_1250 : std_logic_vector(7 downto 0);
    signal conv386_1260 : std_logic_vector(7 downto 0);
    signal conv38_159 : std_logic_vector(15 downto 0);
    signal conv392_1270 : std_logic_vector(7 downto 0);
    signal conv398_1280 : std_logic_vector(7 downto 0);
    signal conv3_59 : std_logic_vector(15 downto 0);
    signal conv404_1290 : std_logic_vector(7 downto 0);
    signal conv438_1382 : std_logic_vector(7 downto 0);
    signal conv444_1392 : std_logic_vector(7 downto 0);
    signal conv44_171 : std_logic_vector(15 downto 0);
    signal conv450_1402 : std_logic_vector(7 downto 0);
    signal conv456_1412 : std_logic_vector(7 downto 0);
    signal conv462_1422 : std_logic_vector(7 downto 0);
    signal conv468_1432 : std_logic_vector(7 downto 0);
    signal conv474_1442 : std_logic_vector(7 downto 0);
    signal conv47_184 : std_logic_vector(15 downto 0);
    signal conv480_1452 : std_logic_vector(7 downto 0);
    signal conv53_196 : std_logic_vector(15 downto 0);
    signal conv56_209 : std_logic_vector(15 downto 0);
    signal conv61_218 : std_logic_vector(31 downto 0);
    signal conv63_222 : std_logic_vector(31 downto 0);
    signal conv65_226 : std_logic_vector(31 downto 0);
    signal conv82_263 : std_logic_vector(31 downto 0);
    signal conv84_267 : std_logic_vector(31 downto 0);
    signal conv87_271 : std_logic_vector(31 downto 0);
    signal conv8_71 : std_logic_vector(15 downto 0);
    signal conv90_275 : std_logic_vector(31 downto 0);
    signal conv95_297 : std_logic_vector(15 downto 0);
    signal conv98_310 : std_logic_vector(15 downto 0);
    signal exitcond1_1487 : std_logic_vector(0 downto 0);
    signal exitcond2_844 : std_logic_vector(0 downto 0);
    signal exitcond3_637 : std_logic_vector(0 downto 0);
    signal exitcond_956 : std_logic_vector(0 downto 0);
    signal iNsTr_14_248 : std_logic_vector(31 downto 0);
    signal iNsTr_198_1344 : std_logic_vector(63 downto 0);
    signal iNsTr_26_459 : std_logic_vector(63 downto 0);
    signal iNsTr_39_666 : std_logic_vector(63 downto 0);
    signal iNsTr_53_910 : std_logic_vector(63 downto 0);
    signal indvar526_926 : std_logic_vector(63 downto 0);
    signal indvar540_682 : std_logic_vector(63 downto 0);
    signal indvar556_475 : std_logic_vector(63 downto 0);
    signal indvar_1360 : std_logic_vector(63 downto 0);
    signal indvarx_xnext527_951 : std_logic_vector(63 downto 0);
    signal indvarx_xnext541_839 : std_logic_vector(63 downto 0);
    signal indvarx_xnext557_632 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1482 : std_logic_vector(63 downto 0);
    signal mul256_870 : std_logic_vector(31 downto 0);
    signal mul259_875 : std_logic_vector(31 downto 0);
    signal mul66_236 : std_logic_vector(31 downto 0);
    signal mul85_280 : std_logic_vector(31 downto 0);
    signal mul88_285 : std_logic_vector(31 downto 0);
    signal mul91_290 : std_logic_vector(31 downto 0);
    signal mul_231 : std_logic_vector(31 downto 0);
    signal ptr_deref_1377_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1377_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1377_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1377_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1377_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_624_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_624_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_624_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_624_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_624_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_624_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_831_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_831_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_831_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_831_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_831_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_831_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_942_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_942_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_942_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_942_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_942_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_942_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_328 : std_logic_vector(15 downto 0);
    signal shl114_353 : std_logic_vector(15 downto 0);
    signal shl123_378 : std_logic_vector(15 downto 0);
    signal shl132_403 : std_logic_vector(15 downto 0);
    signal shl146_502 : std_logic_vector(63 downto 0);
    signal shl152_520 : std_logic_vector(63 downto 0);
    signal shl158_538 : std_logic_vector(63 downto 0);
    signal shl164_556 : std_logic_vector(63 downto 0);
    signal shl170_574 : std_logic_vector(63 downto 0);
    signal shl176_592 : std_logic_vector(63 downto 0);
    signal shl182_610 : std_logic_vector(63 downto 0);
    signal shl18_102 : std_logic_vector(15 downto 0);
    signal shl202_709 : std_logic_vector(63 downto 0);
    signal shl208_727 : std_logic_vector(63 downto 0);
    signal shl214_745 : std_logic_vector(63 downto 0);
    signal shl220_763 : std_logic_vector(63 downto 0);
    signal shl226_781 : std_logic_vector(63 downto 0);
    signal shl232_799 : std_logic_vector(63 downto 0);
    signal shl238_817 : std_logic_vector(63 downto 0);
    signal shl27_127 : std_logic_vector(15 downto 0);
    signal shl36_152 : std_logic_vector(15 downto 0);
    signal shl45_177 : std_logic_vector(15 downto 0);
    signal shl54_202 : std_logic_vector(15 downto 0);
    signal shl96_303 : std_logic_vector(15 downto 0);
    signal shl9_77 : std_logic_vector(15 downto 0);
    signal shl_52 : std_logic_vector(15 downto 0);
    signal shr304_1052 : std_logic_vector(31 downto 0);
    signal shr321_1108 : std_logic_vector(31 downto 0);
    signal shr338_1164 : std_logic_vector(31 downto 0);
    signal shr365_1226 : std_logic_vector(63 downto 0);
    signal shr371_1236 : std_logic_vector(63 downto 0);
    signal shr377_1246 : std_logic_vector(63 downto 0);
    signal shr383_1256 : std_logic_vector(63 downto 0);
    signal shr389_1266 : std_logic_vector(63 downto 0);
    signal shr395_1276 : std_logic_vector(63 downto 0);
    signal shr401_1286 : std_logic_vector(63 downto 0);
    signal shr441_1388 : std_logic_vector(63 downto 0);
    signal shr447_1398 : std_logic_vector(63 downto 0);
    signal shr453_1408 : std_logic_vector(63 downto 0);
    signal shr459_1418 : std_logic_vector(63 downto 0);
    signal shr465_1428 : std_logic_vector(63 downto 0);
    signal shr471_1438 : std_logic_vector(63 downto 0);
    signal shr477_1448 : std_logic_vector(63 downto 0);
    signal shr_242 : std_logic_vector(31 downto 0);
    signal sub_1213 : std_logic_vector(63 downto 0);
    signal tmp434_1378 : std_logic_vector(63 downto 0);
    signal tmp521_1328 : std_logic_vector(31 downto 0);
    signal tmp521x_xop_1340 : std_logic_vector(31 downto 0);
    signal tmp522_1334 : std_logic_vector(0 downto 0);
    signal tmp525_1357 : std_logic_vector(63 downto 0);
    signal tmp533_894 : std_logic_vector(31 downto 0);
    signal tmp533x_xop_906 : std_logic_vector(31 downto 0);
    signal tmp534_900 : std_logic_vector(0 downto 0);
    signal tmp538_923 : std_logic_vector(63 downto 0);
    signal tmp549_650 : std_logic_vector(31 downto 0);
    signal tmp549x_xop_662 : std_logic_vector(31 downto 0);
    signal tmp550_656 : std_logic_vector(0 downto 0);
    signal tmp554_679 : std_logic_vector(63 downto 0);
    signal tmp563x_xop_455 : std_logic_vector(31 downto 0);
    signal tmp564_449 : std_logic_vector(0 downto 0);
    signal tmp568_472 : std_logic_vector(63 downto 0);
    signal type_cast_1005_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1009_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_100_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1050_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1162_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1206_wire : std_logic_vector(63 downto 0);
    signal type_cast_1224_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1234_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1244_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_125_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1264_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1274_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1284_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1332_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1348_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1355_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1364_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1366_wire : std_logic_vector(63 downto 0);
    signal type_cast_1386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1396_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1416_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1426_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1480_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_150_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_175_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_200_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_240_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_252_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_301_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_326_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_351_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_376_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_401_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_434_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_453_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_470_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_479_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_481_wire : std_logic_vector(63 downto 0);
    signal type_cast_500_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_50_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_536_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_554_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_572_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_590_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_630_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_670_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_677_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_685_wire : std_logic_vector(63 downto 0);
    signal type_cast_688_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_707_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_725_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_743_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_75_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_761_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_779_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_797_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_815_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_837_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_879_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_904_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_914_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_921_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_929_wire : std_logic_vector(63 downto 0);
    signal type_cast_932_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_949_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_972_wire : std_logic_vector(63 downto 0);
    signal xx_xop570_916 : std_logic_vector(63 downto 0);
    signal xx_xop571_672 : std_logic_vector(63 downto 0);
    signal xx_xop572_465 : std_logic_vector(63 downto 0);
    signal xx_xop_1350 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1372_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1372_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1372_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1372_resized_base_address <= "00000000000000";
    array_obj_ref_487_constant_part_of_offset <= "00000000000000";
    array_obj_ref_487_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_487_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_487_resized_base_address <= "00000000000000";
    array_obj_ref_694_constant_part_of_offset <= "00000100010";
    array_obj_ref_694_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_694_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_694_resized_base_address <= "00000000000";
    array_obj_ref_938_constant_part_of_offset <= "00000000000000";
    array_obj_ref_938_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_938_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_938_resized_base_address <= "00000000000000";
    ptr_deref_1377_word_offset_0 <= "00000000000000";
    ptr_deref_624_word_offset_0 <= "00000000000000";
    ptr_deref_831_word_offset_0 <= "00000000000";
    ptr_deref_942_word_offset_0 <= "00000000000000";
    type_cast_1005_wire_constant <= "0000000000000000";
    type_cast_1009_wire_constant <= "0000000000000000";
    type_cast_100_wire_constant <= "0000000000001000";
    type_cast_1050_wire_constant <= "00000000000000000000000000010010";
    type_cast_1106_wire_constant <= "00000000000000000000000000010001";
    type_cast_1162_wire_constant <= "00000000000000000000000000010000";
    type_cast_1224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1234_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1244_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1254_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_125_wire_constant <= "0000000000001000";
    type_cast_1264_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1274_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1284_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1326_wire_constant <= "00000000000000000000000000000010";
    type_cast_1332_wire_constant <= "00000000000000000000000000000001";
    type_cast_1338_wire_constant <= "11111111111111111111111111111111";
    type_cast_1348_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1355_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1406_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1416_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1426_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1446_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1480_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_150_wire_constant <= "0000000000001000";
    type_cast_175_wire_constant <= "0000000000001000";
    type_cast_200_wire_constant <= "0000000000001000";
    type_cast_240_wire_constant <= "00000000000000000000000000000010";
    type_cast_246_wire_constant <= "00000000000000000000000000000001";
    type_cast_252_wire_constant <= "01111111111111111111111111111110";
    type_cast_301_wire_constant <= "0000000000001000";
    type_cast_326_wire_constant <= "0000000000001000";
    type_cast_351_wire_constant <= "0000000000001000";
    type_cast_376_wire_constant <= "0000000000001000";
    type_cast_401_wire_constant <= "0000000000001000";
    type_cast_419_wire_constant <= "00000000000000000000000000000011";
    type_cast_434_wire_constant <= "00000000000000000000000000000011";
    type_cast_447_wire_constant <= "00000000000000000000000000000001";
    type_cast_453_wire_constant <= "11111111111111111111111111111111";
    type_cast_463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_470_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_479_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_500_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_50_wire_constant <= "0000000000001000";
    type_cast_518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_536_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_554_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_572_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_590_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_630_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_648_wire_constant <= "00000000000000000000000000000010";
    type_cast_654_wire_constant <= "00000000000000000000000000000001";
    type_cast_660_wire_constant <= "11111111111111111111111111111111";
    type_cast_670_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_677_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_688_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_707_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_725_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_743_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_75_wire_constant <= "0000000000001000";
    type_cast_761_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_779_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_797_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_815_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_837_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_879_wire_constant <= "00000000000000000000000000000011";
    type_cast_892_wire_constant <= "00000000000000000000000000000010";
    type_cast_898_wire_constant <= "00000000000000000000000000000001";
    type_cast_904_wire_constant <= "11111111111111111111111111111111";
    type_cast_914_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_921_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_932_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_944_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_949_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1360: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1364_wire_constant & type_cast_1366_wire;
      req <= phi_stmt_1360_req_0 & phi_stmt_1360_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1360",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1360_ack_0,
          idata => idata,
          odata => indvar_1360,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1360
    phi_stmt_475: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_479_wire_constant & type_cast_481_wire;
      req <= phi_stmt_475_req_0 & phi_stmt_475_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_475",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_475_ack_0,
          idata => idata,
          odata => indvar556_475,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_475
    phi_stmt_682: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_685_wire & type_cast_688_wire_constant;
      req <= phi_stmt_682_req_0 & phi_stmt_682_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_682",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_682_ack_0,
          idata => idata,
          odata => indvar540_682,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_682
    phi_stmt_926: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_929_wire & type_cast_932_wire_constant;
      req <= phi_stmt_926_req_0 & phi_stmt_926_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_926",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_926_ack_0,
          idata => idata,
          odata => indvar526_926,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_926
    -- flow-through select operator MUX_1356_inst
    tmp525_1357 <= xx_xop_1350 when (tmp522_1334(0) /=  '0') else type_cast_1355_wire_constant;
    -- flow-through select operator MUX_471_inst
    tmp568_472 <= xx_xop572_465 when (tmp564_449(0) /=  '0') else type_cast_470_wire_constant;
    -- flow-through select operator MUX_678_inst
    tmp554_679 <= xx_xop571_672 when (tmp550_656(0) /=  '0') else type_cast_677_wire_constant;
    -- flow-through select operator MUX_922_inst
    tmp538_923 <= xx_xop570_916 when (tmp534_900(0) /=  '0') else type_cast_921_wire_constant;
    addr_of_1373_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1373_final_reg_req_0;
      addr_of_1373_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1373_final_reg_req_1;
      addr_of_1373_final_reg_ack_1<= rack(0);
      addr_of_1373_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1373_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1372_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx433_1374,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_488_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_488_final_reg_req_0;
      addr_of_488_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_488_final_reg_req_1;
      addr_of_488_final_reg_ack_1<= rack(0);
      addr_of_488_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_488_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_487_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_695_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_695_final_reg_req_0;
      addr_of_695_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_695_final_reg_req_1;
      addr_of_695_final_reg_ack_1<= rack(0);
      addr_of_695_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_695_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_694_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_939_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_939_final_reg_req_0;
      addr_of_939_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_939_final_reg_req_1;
      addr_of_939_final_reg_ack_1<= rack(0);
      addr_of_939_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_939_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_938_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_940,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1062_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1062_inst_req_0;
      type_cast_1062_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1062_inst_req_1;
      type_cast_1062_inst_ack_1<= rack(0);
      type_cast_1062_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1062_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_242,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1063,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_108_inst_req_0;
      type_cast_108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_108_inst_req_1;
      type_cast_108_inst_ack_1<= rack(0);
      type_cast_108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1111_inst_req_0;
      type_cast_1111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1111_inst_req_1;
      type_cast_1111_inst_ack_1<= rack(0);
      type_cast_1111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1118_inst_req_0;
      type_cast_1118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1118_inst_req_1;
      type_cast_1118_inst_ack_1<= rack(0);
      type_cast_1118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1164,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1174_inst_req_0;
      type_cast_1174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1174_inst_req_1;
      type_cast_1174_inst_ack_1<= rack(0);
      type_cast_1174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1207_inst_req_0;
      type_cast_1207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1207_inst_req_1;
      type_cast_1207_inst_ack_1<= rack(0);
      type_cast_1207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1206_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_120_inst_req_0;
      type_cast_120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_120_inst_req_1;
      type_cast_120_inst_ack_1<= rack(0);
      type_cast_120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1219_inst_req_0;
      type_cast_1219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1219_inst_req_1;
      type_cast_1219_inst_ack_1<= rack(0);
      type_cast_1219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv362_1220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1229_inst_req_0;
      type_cast_1229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1229_inst_req_1;
      type_cast_1229_inst_ack_1<= rack(0);
      type_cast_1229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr365_1226,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv368_1230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1239_inst_req_0;
      type_cast_1239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1239_inst_req_1;
      type_cast_1239_inst_ack_1<= rack(0);
      type_cast_1239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr371_1236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv374_1240,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1249_inst_req_0;
      type_cast_1249_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1249_inst_req_1;
      type_cast_1249_inst_ack_1<= rack(0);
      type_cast_1249_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr377_1246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv380_1250,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1259_inst_req_0;
      type_cast_1259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1259_inst_req_1;
      type_cast_1259_inst_ack_1<= rack(0);
      type_cast_1259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr383_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv386_1260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1269_inst_req_0;
      type_cast_1269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1269_inst_req_1;
      type_cast_1269_inst_ack_1<= rack(0);
      type_cast_1269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr389_1266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv392_1270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr395_1276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv398_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1289_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1289_inst_req_0;
      type_cast_1289_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1289_inst_req_1;
      type_cast_1289_inst_ack_1<= rack(0);
      type_cast_1289_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1289_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr401_1286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv404_1290,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_133_inst_req_0;
      type_cast_133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_133_inst_req_1;
      type_cast_133_inst_ack_1<= rack(0);
      type_cast_133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_133_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1343_inst_req_0;
      type_cast_1343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1343_inst_req_1;
      type_cast_1343_inst_ack_1<= rack(0);
      type_cast_1343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp521x_xop_1340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_198_1344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1366_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1381_inst_req_0;
      type_cast_1381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1381_inst_req_1;
      type_cast_1381_inst_ack_1<= rack(0);
      type_cast_1381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp434_1378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv438_1382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1391_inst_req_0;
      type_cast_1391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1391_inst_req_1;
      type_cast_1391_inst_ack_1<= rack(0);
      type_cast_1391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr441_1388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv444_1392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1401_inst_req_0;
      type_cast_1401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1401_inst_req_1;
      type_cast_1401_inst_ack_1<= rack(0);
      type_cast_1401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr447_1398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv450_1402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1411_inst_req_0;
      type_cast_1411_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1411_inst_req_1;
      type_cast_1411_inst_ack_1<= rack(0);
      type_cast_1411_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1411_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr453_1408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv456_1412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1421_inst_req_0;
      type_cast_1421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1421_inst_req_1;
      type_cast_1421_inst_ack_1<= rack(0);
      type_cast_1421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr459_1418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv462_1422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1431_inst_req_0;
      type_cast_1431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1431_inst_req_1;
      type_cast_1431_inst_ack_1<= rack(0);
      type_cast_1431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr465_1428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv468_1432,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1441_inst_req_0;
      type_cast_1441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1441_inst_req_1;
      type_cast_1441_inst_ack_1<= rack(0);
      type_cast_1441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr471_1438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv474_1442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1451_inst_req_0;
      type_cast_1451_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1451_inst_req_1;
      type_cast_1451_inst_ack_1<= rack(0);
      type_cast_1451_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1451_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr477_1448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv480_1452,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_145_inst_req_0;
      type_cast_145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_145_inst_req_1;
      type_cast_145_inst_ack_1<= rack(0);
      type_cast_145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_158_inst_req_0;
      type_cast_158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_158_inst_req_1;
      type_cast_158_inst_ack_1<= rack(0);
      type_cast_158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_170_inst_req_0;
      type_cast_170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_170_inst_req_1;
      type_cast_170_inst_ack_1<= rack(0);
      type_cast_170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_183_inst_req_0;
      type_cast_183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_183_inst_req_1;
      type_cast_183_inst_ack_1<= rack(0);
      type_cast_183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_195_inst_req_0;
      type_cast_195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_195_inst_req_1;
      type_cast_195_inst_ack_1<= rack(0);
      type_cast_195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_208_inst_req_0;
      type_cast_208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_208_inst_req_1;
      type_cast_208_inst_ack_1<= rack(0);
      type_cast_208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_217_inst_req_0;
      type_cast_217_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_217_inst_req_1;
      type_cast_217_inst_ack_1<= rack(0);
      type_cast_217_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_217_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_64,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_221_inst_req_0;
      type_cast_221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_221_inst_req_1;
      type_cast_221_inst_ack_1<= rack(0);
      type_cast_221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_89,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_225_inst_req_0;
      type_cast_225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_225_inst_req_1;
      type_cast_225_inst_ack_1<= rack(0);
      type_cast_225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_262_inst_req_0;
      type_cast_262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_262_inst_req_1;
      type_cast_262_inst_ack_1<= rack(0);
      type_cast_262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_139,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_266_inst_req_0;
      type_cast_266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_266_inst_req_1;
      type_cast_266_inst_ack_1<= rack(0);
      type_cast_266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_164,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_270_inst_req_0;
      type_cast_270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_270_inst_req_1;
      type_cast_270_inst_ack_1<= rack(0);
      type_cast_270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_274_inst_req_0;
      type_cast_274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_274_inst_req_1;
      type_cast_274_inst_ack_1<= rack(0);
      type_cast_274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_296_inst_req_0;
      type_cast_296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_296_inst_req_1;
      type_cast_296_inst_ack_1<= rack(0);
      type_cast_296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_296_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_309_inst_req_0;
      type_cast_309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_309_inst_req_1;
      type_cast_309_inst_ack_1<= rack(0);
      type_cast_309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_321_inst_req_0;
      type_cast_321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_321_inst_req_1;
      type_cast_321_inst_ack_1<= rack(0);
      type_cast_321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_334_inst_req_0;
      type_cast_334_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_334_inst_req_1;
      type_cast_334_inst_ack_1<= rack(0);
      type_cast_334_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_334_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_331,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_346_inst_req_0;
      type_cast_346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_346_inst_req_1;
      type_cast_346_inst_ack_1<= rack(0);
      type_cast_346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_359_inst_req_0;
      type_cast_359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_359_inst_req_1;
      type_cast_359_inst_ack_1<= rack(0);
      type_cast_359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_384_inst_req_0;
      type_cast_384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_384_inst_req_1;
      type_cast_384_inst_ack_1<= rack(0);
      type_cast_384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_396_inst_req_0;
      type_cast_396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_396_inst_req_1;
      type_cast_396_inst_ack_1<= rack(0);
      type_cast_396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_409_inst_req_0;
      type_cast_409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_409_inst_req_1;
      type_cast_409_inst_ack_1<= rack(0);
      type_cast_409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_458_inst_req_0;
      type_cast_458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_458_inst_req_1;
      type_cast_458_inst_ack_1<= rack(0);
      type_cast_458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp563x_xop_455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_459,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_45_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_45_inst_req_0;
      type_cast_45_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_45_inst_req_1;
      type_cast_45_inst_ack_1<= rack(0);
      type_cast_45_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_45_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_42,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_46,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_481_inst_req_0;
      type_cast_481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_481_inst_req_1;
      type_cast_481_inst_ack_1<= rack(0);
      type_cast_481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext557_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_481_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_495_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_495_inst_req_0;
      type_cast_495_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_495_inst_req_1;
      type_cast_495_inst_ack_1<= rack(0);
      type_cast_495_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_495_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_496,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_508_inst_req_0;
      type_cast_508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_508_inst_req_1;
      type_cast_508_inst_ack_1<= rack(0);
      type_cast_508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_526_inst_req_0;
      type_cast_526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_526_inst_req_1;
      type_cast_526_inst_ack_1<= rack(0);
      type_cast_526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_526_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_527,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_544_inst_req_0;
      type_cast_544_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_544_inst_req_1;
      type_cast_544_inst_ack_1<= rack(0);
      type_cast_544_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_544_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_562_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_562_inst_req_0;
      type_cast_562_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_562_inst_req_1;
      type_cast_562_inst_ack_1<= rack(0);
      type_cast_562_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_562_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_559,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_563,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_580_inst_req_0;
      type_cast_580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_580_inst_req_1;
      type_cast_580_inst_ack_1<= rack(0);
      type_cast_580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_58_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_58_inst_req_0;
      type_cast_58_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_58_inst_req_1;
      type_cast_58_inst_ack_1<= rack(0);
      type_cast_58_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_58_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_55,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_59,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_598_inst_req_0;
      type_cast_598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_598_inst_req_1;
      type_cast_598_inst_ack_1<= rack(0);
      type_cast_598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_616_inst_req_0;
      type_cast_616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_616_inst_req_1;
      type_cast_616_inst_ack_1<= rack(0);
      type_cast_616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_665_inst_req_0;
      type_cast_665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_665_inst_req_1;
      type_cast_665_inst_ack_1<= rack(0);
      type_cast_665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp549x_xop_662,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_685_inst_req_0;
      type_cast_685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_685_inst_req_1;
      type_cast_685_inst_ack_1<= rack(0);
      type_cast_685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext541_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_685_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_702_inst_req_0;
      type_cast_702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_702_inst_req_1;
      type_cast_702_inst_ack_1<= rack(0);
      type_cast_702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_70_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_70_inst_req_0;
      type_cast_70_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_70_inst_req_1;
      type_cast_70_inst_ack_1<= rack(0);
      type_cast_70_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_70_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_71,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_715_inst_req_0;
      type_cast_715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_715_inst_req_1;
      type_cast_715_inst_ack_1<= rack(0);
      type_cast_715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_712,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_733_inst_req_0;
      type_cast_733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_733_inst_req_1;
      type_cast_733_inst_ack_1<= rack(0);
      type_cast_733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_769_inst_req_0;
      type_cast_769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_769_inst_req_1;
      type_cast_769_inst_ack_1<= rack(0);
      type_cast_769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_766,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_787_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_787_inst_req_0;
      type_cast_787_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_787_inst_req_1;
      type_cast_787_inst_ack_1<= rack(0);
      type_cast_787_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_787_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_784,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_805_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_805_inst_req_0;
      type_cast_805_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_805_inst_req_1;
      type_cast_805_inst_ack_1<= rack(0);
      type_cast_805_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_805_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_802,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_806,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_823_inst_req_0;
      type_cast_823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_823_inst_req_1;
      type_cast_823_inst_ack_1<= rack(0);
      type_cast_823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_80,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_84,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_856_inst_req_0;
      type_cast_856_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_856_inst_req_1;
      type_cast_856_inst_ack_1<= rack(0);
      type_cast_856_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_856_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_857,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_860_inst_req_0;
      type_cast_860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_860_inst_req_1;
      type_cast_860_inst_ack_1<= rack(0);
      type_cast_860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_861,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_864_inst_req_0;
      type_cast_864_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_864_inst_req_1;
      type_cast_864_inst_ack_1<= rack(0);
      type_cast_864_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_865,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_909_inst_req_0;
      type_cast_909_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_909_inst_req_1;
      type_cast_909_inst_ack_1<= rack(0);
      type_cast_909_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp533x_xop_906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_910,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_929_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_929_inst_req_0;
      type_cast_929_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_929_inst_req_1;
      type_cast_929_inst_ack_1<= rack(0);
      type_cast_929_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_929_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext527_951,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_929_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_973_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_973_inst_req_0;
      type_cast_973_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_973_inst_req_1;
      type_cast_973_inst_ack_1<= rack(0);
      type_cast_973_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_973_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_972_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_974,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1372_index_1_rename
    process(R_indvar_1371_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1371_resized;
      ov(13 downto 0) := iv;
      R_indvar_1371_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1372_index_1_resize
    process(indvar_1360) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1360;
      ov := iv(13 downto 0);
      R_indvar_1371_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1372_root_address_inst
    process(array_obj_ref_1372_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1372_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1372_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_487_index_1_rename
    process(R_indvar556_486_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar556_486_resized;
      ov(13 downto 0) := iv;
      R_indvar556_486_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_487_index_1_resize
    process(indvar556_475) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar556_475;
      ov := iv(13 downto 0);
      R_indvar556_486_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_487_root_address_inst
    process(array_obj_ref_487_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_487_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_487_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_694_index_1_rename
    process(R_indvar540_693_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar540_693_resized;
      ov(10 downto 0) := iv;
      R_indvar540_693_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_694_index_1_resize
    process(indvar540_682) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar540_682;
      ov := iv(10 downto 0);
      R_indvar540_693_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_694_root_address_inst
    process(array_obj_ref_694_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_694_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_694_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_938_index_1_rename
    process(R_indvar526_937_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar526_937_resized;
      ov(13 downto 0) := iv;
      R_indvar526_937_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_938_index_1_resize
    process(indvar526_926) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar526_926;
      ov := iv(13 downto 0);
      R_indvar526_937_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_938_root_address_inst
    process(array_obj_ref_938_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_938_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_938_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1377_addr_0
    process(ptr_deref_1377_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1377_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1377_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1377_base_resize
    process(arrayidx433_1374) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx433_1374;
      ov := iv(13 downto 0);
      ptr_deref_1377_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1377_gather_scatter
    process(ptr_deref_1377_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1377_data_0;
      ov(63 downto 0) := iv;
      tmp434_1378 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1377_root_address_inst
    process(ptr_deref_1377_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1377_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1377_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_addr_0
    process(ptr_deref_624_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_624_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_624_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_base_resize
    process(arrayidx_489) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_489;
      ov := iv(13 downto 0);
      ptr_deref_624_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_gather_scatter
    process(add186_622) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_622;
      ov(63 downto 0) := iv;
      ptr_deref_624_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_624_root_address_inst
    process(ptr_deref_624_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_624_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_624_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_addr_0
    process(ptr_deref_831_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_831_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_base_resize
    process(arrayidx246_696) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_696;
      ov := iv(10 downto 0);
      ptr_deref_831_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_gather_scatter
    process(add242_829) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_829;
      ov(63 downto 0) := iv;
      ptr_deref_831_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_root_address_inst
    process(ptr_deref_831_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_831_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_addr_0
    process(ptr_deref_942_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_942_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_base_resize
    process(arrayidx269_940) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_940;
      ov := iv(13 downto 0);
      ptr_deref_942_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_gather_scatter
    process(type_cast_944_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_944_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_942_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_root_address_inst
    process(ptr_deref_942_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_942_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1316_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264506_881;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1316_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1316_branch_req_0,
          ack0 => if_stmt_1316_branch_ack_0,
          ack1 => if_stmt_1316_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1488_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1487;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1488_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1488_branch_req_0,
          ack0 => if_stmt_1488_branch_ack_0,
          ack1 => if_stmt_1488_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_422_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp514_421;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_422_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_422_branch_req_0,
          ack0 => if_stmt_422_branch_ack_0,
          ack1 => if_stmt_422_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_437_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194510_436;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_437_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_437_branch_req_0,
          ack0 => if_stmt_437_branch_ack_0,
          ack1 => if_stmt_437_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_638_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_637;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_638_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_638_branch_req_0,
          ack0 => if_stmt_638_branch_ack_0,
          ack1 => if_stmt_638_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_845_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_844;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_845_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_845_branch_req_0,
          ack0 => if_stmt_845_branch_ack_0,
          ack1 => if_stmt_845_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_882_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264506_881;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_882_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_882_branch_req_0,
          ack0 => if_stmt_882_branch_ack_0,
          ack1 => if_stmt_882_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_957_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_956;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_957_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_957_branch_req_0,
          ack0 => if_stmt_957_branch_ack_0,
          ack1 => if_stmt_957_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1339_inst
    process(tmp521_1328) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp521_1328, type_cast_1338_wire_constant, tmp_var);
      tmp521x_xop_1340 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_258_inst
    process(add74_254, shr_242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_254, shr_242, tmp_var);
      add79_259 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_454_inst
    process(shr_242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_242, type_cast_453_wire_constant, tmp_var);
      tmp563x_xop_455 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_661_inst
    process(tmp549_650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp549_650, type_cast_660_wire_constant, tmp_var);
      tmp549x_xop_662 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_905_inst
    process(tmp533_894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp533_894, type_cast_904_wire_constant, tmp_var);
      tmp533x_xop_906 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1349_inst
    process(iNsTr_198_1344) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_198_1344, type_cast_1348_wire_constant, tmp_var);
      xx_xop_1350 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1481_inst
    process(indvar_1360) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1360, type_cast_1480_wire_constant, tmp_var);
      indvarx_xnext_1482 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_464_inst
    process(iNsTr_26_459) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_459, type_cast_463_wire_constant, tmp_var);
      xx_xop572_465 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_631_inst
    process(indvar556_475) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar556_475, type_cast_630_wire_constant, tmp_var);
      indvarx_xnext557_632 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_671_inst
    process(iNsTr_39_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_666, type_cast_670_wire_constant, tmp_var);
      xx_xop571_672 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_838_inst
    process(indvar540_682) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar540_682, type_cast_837_wire_constant, tmp_var);
      indvarx_xnext541_839 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_915_inst
    process(iNsTr_53_910) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_910, type_cast_914_wire_constant, tmp_var);
      xx_xop570_916 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_950_inst
    process(indvar526_926) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar526_926, type_cast_949_wire_constant, tmp_var);
      indvarx_xnext527_951 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_253_inst
    process(iNsTr_14_248) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_248, type_cast_252_wire_constant, tmp_var);
      add74_254 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1486_inst
    process(indvarx_xnext_1482, tmp525_1357) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1482, tmp525_1357, tmp_var);
      exitcond1_1487 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_636_inst
    process(indvarx_xnext557_632, tmp568_472) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext557_632, tmp568_472, tmp_var);
      exitcond3_637 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_843_inst
    process(indvarx_xnext541_839, tmp554_679) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext541_839, tmp554_679, tmp_var);
      exitcond2_844 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_955_inst
    process(indvarx_xnext527_951, tmp538_923) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext527_951, tmp538_923, tmp_var);
      exitcond_956 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1051_inst
    process(mul66_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_236, type_cast_1050_wire_constant, tmp_var);
      shr304_1052 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1107_inst
    process(mul66_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_236, type_cast_1106_wire_constant, tmp_var);
      shr321_1108 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1163_inst
    process(add79_259) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_259, type_cast_1162_wire_constant, tmp_var);
      shr338_1164 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1327_inst
    process(mul259_875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_875, type_cast_1326_wire_constant, tmp_var);
      tmp521_1328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_241_inst
    process(mul66_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_236, type_cast_240_wire_constant, tmp_var);
      shr_242 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_247_inst
    process(mul66_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_236, type_cast_246_wire_constant, tmp_var);
      iNsTr_14_248 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_649_inst
    process(mul91_290) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_290, type_cast_648_wire_constant, tmp_var);
      tmp549_650 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_893_inst
    process(mul259_875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_875, type_cast_892_wire_constant, tmp_var);
      tmp533_894 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1225_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1224_wire_constant, tmp_var);
      shr365_1226 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1235_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1234_wire_constant, tmp_var);
      shr371_1236 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1245_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1244_wire_constant, tmp_var);
      shr377_1246 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1255_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1254_wire_constant, tmp_var);
      shr383_1256 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1265_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1264_wire_constant, tmp_var);
      shr389_1266 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1275_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1274_wire_constant, tmp_var);
      shr395_1276 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1285_inst
    process(sub_1213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1213, type_cast_1284_wire_constant, tmp_var);
      shr401_1286 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1387_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1386_wire_constant, tmp_var);
      shr441_1388 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1397_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1396_wire_constant, tmp_var);
      shr447_1398 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1407_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1406_wire_constant, tmp_var);
      shr453_1408 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1417_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1416_wire_constant, tmp_var);
      shr459_1418 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1427_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1426_wire_constant, tmp_var);
      shr465_1428 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1437_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1436_wire_constant, tmp_var);
      shr471_1438 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1447_inst
    process(tmp434_1378) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp434_1378, type_cast_1446_wire_constant, tmp_var);
      shr477_1448 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_230_inst
    process(conv63_222, conv61_218) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_222, conv61_218, tmp_var);
      mul_231 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_235_inst
    process(mul_231, conv65_226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_231, conv65_226, tmp_var);
      mul66_236 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_279_inst
    process(conv84_267, conv82_263) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_267, conv82_263, tmp_var);
      mul85_280 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_284_inst
    process(mul85_280, conv87_271) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_280, conv87_271, tmp_var);
      mul88_285 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_289_inst
    process(mul88_285, conv90_275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_285, conv90_275, tmp_var);
      mul91_290 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_869_inst
    process(conv255_861, conv253_857) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_861, conv253_857, tmp_var);
      mul256_870 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_874_inst
    process(mul256_870, conv258_865) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_870, conv258_865, tmp_var);
      mul259_875 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_113_inst
    process(shl18_102, conv20_109) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_102, conv20_109, tmp_var);
      add21_114 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_138_inst
    process(shl27_127, conv29_134) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_127, conv29_134, tmp_var);
      add30_139 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_163_inst
    process(shl36_152, conv38_159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_152, conv38_159, tmp_var);
      add39_164 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_188_inst
    process(shl45_177, conv47_184) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_177, conv47_184, tmp_var);
      add48_189 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_213_inst
    process(shl54_202, conv56_209) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_202, conv56_209, tmp_var);
      add57_214 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_314_inst
    process(shl96_303, conv98_310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_303, conv98_310, tmp_var);
      add99_315 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_339_inst
    process(shl105_328, conv107_335) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_328, conv107_335, tmp_var);
      add108_340 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_364_inst
    process(shl114_353, conv116_360) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_353, conv116_360, tmp_var);
      add117_365 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_389_inst
    process(shl123_378, conv125_385) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_378, conv125_385, tmp_var);
      add126_390 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_414_inst
    process(shl132_403, conv134_410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_403, conv134_410, tmp_var);
      add135_415 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_63_inst
    process(shl_52, conv3_59) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_52, conv3_59, tmp_var);
      add_64 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_88_inst
    process(shl9_77, conv11_84) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_77, conv11_84, tmp_var);
      add12_89 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_513_inst
    process(shl146_502, conv149_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_502, conv149_509, tmp_var);
      add150_514 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_531_inst
    process(shl152_520, conv155_527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_520, conv155_527, tmp_var);
      add156_532 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_549_inst
    process(shl158_538, conv161_545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_538, conv161_545, tmp_var);
      add162_550 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_567_inst
    process(shl164_556, conv167_563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_556, conv167_563, tmp_var);
      add168_568 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_585_inst
    process(shl170_574, conv173_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_574, conv173_581, tmp_var);
      add174_586 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_603_inst
    process(shl176_592, conv179_599) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_592, conv179_599, tmp_var);
      add180_604 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_621_inst
    process(shl182_610, conv185_617) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_610, conv185_617, tmp_var);
      add186_622 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_720_inst
    process(shl202_709, conv205_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_709, conv205_716, tmp_var);
      add206_721 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_738_inst
    process(shl208_727, conv211_734) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_727, conv211_734, tmp_var);
      add212_739 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_756_inst
    process(shl214_745, conv217_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_745, conv217_752, tmp_var);
      add218_757 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_774_inst
    process(shl220_763, conv223_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_763, conv223_770, tmp_var);
      add224_775 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_792_inst
    process(shl226_781, conv229_788) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_781, conv229_788, tmp_var);
      add230_793 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_810_inst
    process(shl232_799, conv235_806) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_799, conv235_806, tmp_var);
      add236_811 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_828_inst
    process(shl238_817, conv241_824) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_817, conv241_824, tmp_var);
      add242_829 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_101_inst
    process(conv17_96) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_96, type_cast_100_wire_constant, tmp_var);
      shl18_102 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_126_inst
    process(conv26_121) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_121, type_cast_125_wire_constant, tmp_var);
      shl27_127 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_151_inst
    process(conv35_146) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_146, type_cast_150_wire_constant, tmp_var);
      shl36_152 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_176_inst
    process(conv44_171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_171, type_cast_175_wire_constant, tmp_var);
      shl45_177 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_201_inst
    process(conv53_196) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_196, type_cast_200_wire_constant, tmp_var);
      shl54_202 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_302_inst
    process(conv95_297) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_297, type_cast_301_wire_constant, tmp_var);
      shl96_303 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_327_inst
    process(conv104_322) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_322, type_cast_326_wire_constant, tmp_var);
      shl105_328 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_352_inst
    process(conv113_347) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_347, type_cast_351_wire_constant, tmp_var);
      shl114_353 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_377_inst
    process(conv122_372) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_372, type_cast_376_wire_constant, tmp_var);
      shl123_378 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_402_inst
    process(conv131_397) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_397, type_cast_401_wire_constant, tmp_var);
      shl132_403 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_51_inst
    process(conv1_46) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_46, type_cast_50_wire_constant, tmp_var);
      shl_52 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_76_inst
    process(conv8_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_71, type_cast_75_wire_constant, tmp_var);
      shl9_77 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_501_inst
    process(conv144_496) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_496, type_cast_500_wire_constant, tmp_var);
      shl146_502 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_519_inst
    process(add150_514) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_514, type_cast_518_wire_constant, tmp_var);
      shl152_520 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_537_inst
    process(add156_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_532, type_cast_536_wire_constant, tmp_var);
      shl158_538 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_555_inst
    process(add162_550) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_550, type_cast_554_wire_constant, tmp_var);
      shl164_556 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_573_inst
    process(add168_568) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_568, type_cast_572_wire_constant, tmp_var);
      shl170_574 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_591_inst
    process(add174_586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_586, type_cast_590_wire_constant, tmp_var);
      shl176_592 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_609_inst
    process(add180_604) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_604, type_cast_608_wire_constant, tmp_var);
      shl182_610 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_708_inst
    process(conv200_703) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_703, type_cast_707_wire_constant, tmp_var);
      shl202_709 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_726_inst
    process(add206_721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_721, type_cast_725_wire_constant, tmp_var);
      shl208_727 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_744_inst
    process(add212_739) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_739, type_cast_743_wire_constant, tmp_var);
      shl214_745 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_762_inst
    process(add218_757) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_757, type_cast_761_wire_constant, tmp_var);
      shl220_763 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_780_inst
    process(add224_775) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_775, type_cast_779_wire_constant, tmp_var);
      shl226_781 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_798_inst
    process(add230_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_793, type_cast_797_wire_constant, tmp_var);
      shl232_799 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_816_inst
    process(add236_811) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_811, type_cast_815_wire_constant, tmp_var);
      shl238_817 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1212_inst
    process(conv355_1208, conv276_974) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1208, conv276_974, tmp_var);
      sub_1213 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1333_inst
    process(tmp521_1328) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp521_1328, type_cast_1332_wire_constant, tmp_var);
      tmp522_1334 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_420_inst
    process(mul66_236) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_236, type_cast_419_wire_constant, tmp_var);
      cmp514_421 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_435_inst
    process(mul91_290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_290, type_cast_434_wire_constant, tmp_var);
      cmp194510_436 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_448_inst
    process(shr_242) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_242, type_cast_447_wire_constant, tmp_var);
      tmp564_449 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_655_inst
    process(tmp549_650) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp549_650, type_cast_654_wire_constant, tmp_var);
      tmp550_656 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_880_inst
    process(mul259_875) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_875, type_cast_879_wire_constant, tmp_var);
      cmp264506_881 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_899_inst
    process(tmp533_894) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp533_894, type_cast_898_wire_constant, tmp_var);
      tmp534_900 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1372_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1371_scaled;
      array_obj_ref_1372_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1372_index_offset_req_0;
      array_obj_ref_1372_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1372_index_offset_req_1;
      array_obj_ref_1372_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_487_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar556_486_scaled;
      array_obj_ref_487_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_487_index_offset_req_0;
      array_obj_ref_487_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_487_index_offset_req_1;
      array_obj_ref_487_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_694_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar540_693_scaled;
      array_obj_ref_694_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_694_index_offset_req_0;
      array_obj_ref_694_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_694_index_offset_req_1;
      array_obj_ref_694_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_938_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar526_937_scaled;
      array_obj_ref_938_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_938_index_offset_req_0;
      array_obj_ref_938_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_938_index_offset_req_1;
      array_obj_ref_938_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1206_inst
    process(call354_1203) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1203, tmp_var);
      type_cast_1206_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_972_inst
    process(call275_968) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_968, tmp_var);
      type_cast_972_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1377_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1377_load_0_req_0;
      ptr_deref_1377_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1377_load_0_req_1;
      ptr_deref_1377_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1377_word_address_0;
      ptr_deref_1377_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_624_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_624_store_0_req_0;
      ptr_deref_624_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_624_store_0_req_1;
      ptr_deref_624_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_624_word_address_0;
      data_in <= ptr_deref_624_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_831_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_831_store_0_req_0;
      ptr_deref_831_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_831_store_0_req_1;
      ptr_deref_831_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_831_word_address_0;
      data_in <= ptr_deref_831_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(10 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_942_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_942_store_0_req_0;
      ptr_deref_942_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_942_store_0_req_1;
      ptr_deref_942_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_942_word_address_0;
      data_in <= ptr_deref_942_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1190_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1190_inst_req_0;
      RPIPE_Block0_done_1190_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1190_inst_req_1;
      RPIPE_Block0_done_1190_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1191 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1193_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1193_inst_req_0;
      RPIPE_Block1_done_1193_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1193_inst_req_1;
      RPIPE_Block1_done_1193_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1194 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1196_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1196_inst_req_0;
      RPIPE_Block2_done_1196_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1196_inst_req_1;
      RPIPE_Block2_done_1196_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1197 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1199_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1199_inst_req_0;
      RPIPE_Block3_done_1199_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1199_inst_req_1;
      RPIPE_Block3_done_1199_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1200 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_141_inst RPIPE_ConvTranspose_input_pipe_504_inst RPIPE_ConvTranspose_input_pipe_54_inst RPIPE_ConvTranspose_input_pipe_801_inst RPIPE_ConvTranspose_input_pipe_491_inst RPIPE_ConvTranspose_input_pipe_594_inst RPIPE_ConvTranspose_input_pipe_41_inst RPIPE_ConvTranspose_input_pipe_91_inst RPIPE_ConvTranspose_input_pipe_558_inst RPIPE_ConvTranspose_input_pipe_612_inst RPIPE_ConvTranspose_input_pipe_522_inst RPIPE_ConvTranspose_input_pipe_116_inst RPIPE_ConvTranspose_input_pipe_729_inst RPIPE_ConvTranspose_input_pipe_576_inst RPIPE_ConvTranspose_input_pipe_79_inst RPIPE_ConvTranspose_input_pipe_104_inst RPIPE_ConvTranspose_input_pipe_698_inst RPIPE_ConvTranspose_input_pipe_540_inst RPIPE_ConvTranspose_input_pipe_783_inst RPIPE_ConvTranspose_input_pipe_747_inst RPIPE_ConvTranspose_input_pipe_66_inst RPIPE_ConvTranspose_input_pipe_711_inst RPIPE_ConvTranspose_input_pipe_819_inst RPIPE_ConvTranspose_input_pipe_765_inst RPIPE_ConvTranspose_input_pipe_129_inst RPIPE_ConvTranspose_input_pipe_154_inst RPIPE_ConvTranspose_input_pipe_166_inst RPIPE_ConvTranspose_input_pipe_179_inst RPIPE_ConvTranspose_input_pipe_191_inst RPIPE_ConvTranspose_input_pipe_204_inst RPIPE_ConvTranspose_input_pipe_292_inst RPIPE_ConvTranspose_input_pipe_305_inst RPIPE_ConvTranspose_input_pipe_317_inst RPIPE_ConvTranspose_input_pipe_330_inst RPIPE_ConvTranspose_input_pipe_342_inst RPIPE_ConvTranspose_input_pipe_355_inst RPIPE_ConvTranspose_input_pipe_367_inst RPIPE_ConvTranspose_input_pipe_380_inst RPIPE_ConvTranspose_input_pipe_392_inst RPIPE_ConvTranspose_input_pipe_405_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_504_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_54_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_801_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_491_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_594_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_41_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_558_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_612_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_522_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_729_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_576_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_79_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_104_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_698_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_540_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_783_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_747_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_711_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_819_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_765_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_129_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_154_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_179_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_191_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_204_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_292_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_305_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_317_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_330_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_342_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_355_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_367_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_380_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_392_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_405_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_504_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_54_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_801_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_491_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_594_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_41_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_558_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_612_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_522_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_729_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_576_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_79_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_104_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_698_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_540_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_783_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_747_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_711_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_819_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_765_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_129_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_154_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_179_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_191_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_204_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_292_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_305_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_317_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_330_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_342_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_355_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_367_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_380_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_392_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_405_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_504_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_54_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_801_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_491_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_594_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_41_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_558_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_612_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_522_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_729_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_576_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_79_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_104_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_698_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_540_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_783_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_747_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_711_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_819_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_765_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_129_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_154_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_179_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_191_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_204_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_292_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_305_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_317_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_330_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_342_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_355_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_367_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_380_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_392_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_405_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_504_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_54_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_801_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_491_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_594_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_41_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_558_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_612_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_522_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_729_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_576_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_79_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_104_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_698_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_540_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_783_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_747_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_711_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_819_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_765_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_129_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_154_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_179_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_191_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_204_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_292_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_305_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_317_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_330_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_342_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_355_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_367_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_380_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_392_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_405_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call32_142 <= data_out(319 downto 312);
      call147_505 <= data_out(311 downto 304);
      call2_55 <= data_out(303 downto 296);
      call233_802 <= data_out(295 downto 288);
      call143_492 <= data_out(287 downto 280);
      call177_595 <= data_out(279 downto 272);
      call_42 <= data_out(271 downto 264);
      call14_92 <= data_out(263 downto 256);
      call165_559 <= data_out(255 downto 248);
      call183_613 <= data_out(247 downto 240);
      call153_523 <= data_out(239 downto 232);
      call23_117 <= data_out(231 downto 224);
      call209_730 <= data_out(223 downto 216);
      call171_577 <= data_out(215 downto 208);
      call10_80 <= data_out(207 downto 200);
      call19_105 <= data_out(199 downto 192);
      call199_699 <= data_out(191 downto 184);
      call159_541 <= data_out(183 downto 176);
      call227_784 <= data_out(175 downto 168);
      call215_748 <= data_out(167 downto 160);
      call5_67 <= data_out(159 downto 152);
      call203_712 <= data_out(151 downto 144);
      call239_820 <= data_out(143 downto 136);
      call221_766 <= data_out(135 downto 128);
      call28_130 <= data_out(127 downto 120);
      call37_155 <= data_out(119 downto 112);
      call41_167 <= data_out(111 downto 104);
      call46_180 <= data_out(103 downto 96);
      call50_192 <= data_out(95 downto 88);
      call55_205 <= data_out(87 downto 80);
      call92_293 <= data_out(79 downto 72);
      call97_306 <= data_out(71 downto 64);
      call101_318 <= data_out(63 downto 56);
      call106_331 <= data_out(55 downto 48);
      call110_343 <= data_out(47 downto 40);
      call115_356 <= data_out(39 downto 32);
      call119_368 <= data_out(31 downto 24);
      call124_381 <= data_out(23 downto 16);
      call128_393 <= data_out(15 downto 8);
      call133_406 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_982_inst WPIPE_Block0_start_985_inst WPIPE_Block0_start_988_inst WPIPE_Block0_start_991_inst WPIPE_Block0_start_994_inst WPIPE_Block0_start_1003_inst WPIPE_Block0_start_1007_inst WPIPE_Block0_start_1017_inst WPIPE_Block0_start_997_inst WPIPE_Block0_start_976_inst WPIPE_Block0_start_1000_inst WPIPE_Block0_start_979_inst WPIPE_Block0_start_1014_inst WPIPE_Block0_start_1011_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_982_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_985_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_988_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_991_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_994_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_1003_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_1007_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_1017_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_997_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_976_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_1000_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_979_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_1014_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1011_inst_req_0;
      WPIPE_Block0_start_982_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_985_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_988_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_991_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_994_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_1003_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_1007_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_1017_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_997_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_976_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_1000_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_979_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_1014_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1011_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_982_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_985_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_988_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_991_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_994_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_1003_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_1007_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_1017_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_997_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_976_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_1000_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_979_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_1014_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1011_inst_req_1;
      WPIPE_Block0_start_982_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_985_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_988_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_991_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_994_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_1003_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_1007_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_1017_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_997_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_976_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_1000_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_979_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_1014_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1011_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add21_114 & add30_139 & add39_164 & add48_189 & add57_214 & type_cast_1005_wire_constant & type_cast_1009_wire_constant & add135_415 & add99_315 & add_64 & add108_340 & add12_89 & add126_390 & add117_365;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1020_inst WPIPE_Block1_start_1023_inst WPIPE_Block1_start_1026_inst WPIPE_Block1_start_1038_inst WPIPE_Block1_start_1032_inst WPIPE_Block1_start_1067_inst WPIPE_Block1_start_1064_inst WPIPE_Block1_start_1041_inst WPIPE_Block1_start_1070_inst WPIPE_Block1_start_1035_inst WPIPE_Block1_start_1073_inst WPIPE_Block1_start_1044_inst WPIPE_Block1_start_1029_inst WPIPE_Block1_start_1057_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1020_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1023_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1026_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1038_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1032_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1067_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1064_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1041_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1070_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1035_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1073_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1044_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1029_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1057_inst_req_0;
      WPIPE_Block1_start_1020_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1023_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1026_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1038_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1032_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1067_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1064_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1041_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1070_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1035_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1073_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1044_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1029_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1057_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1020_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1023_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1026_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1038_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1032_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1067_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1064_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1041_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1070_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1035_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1073_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1044_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1029_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1057_inst_req_1;
      WPIPE_Block1_start_1020_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1023_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1026_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1038_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1032_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1067_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1064_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1041_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1070_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1035_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1073_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1044_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1029_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1057_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_64 & add12_89 & add21_114 & add57_214 & add39_164 & add117_365 & conv307_1063 & add99_315 & add126_390 & add48_189 & add135_415 & add108_340 & add30_139 & conv305_1056;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1094_inst WPIPE_Block2_start_1113_inst WPIPE_Block2_start_1123_inst WPIPE_Block2_start_1126_inst WPIPE_Block2_start_1085_inst WPIPE_Block2_start_1091_inst WPIPE_Block2_start_1129_inst WPIPE_Block2_start_1097_inst WPIPE_Block2_start_1100_inst WPIPE_Block2_start_1082_inst WPIPE_Block2_start_1120_inst WPIPE_Block2_start_1088_inst WPIPE_Block2_start_1079_inst WPIPE_Block2_start_1076_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1094_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1113_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1123_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1126_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1085_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1091_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1129_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1097_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1100_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1082_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1120_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1088_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1079_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1076_inst_req_0;
      WPIPE_Block2_start_1094_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1113_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1123_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1126_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1085_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1091_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1129_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1097_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1100_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1082_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1120_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1088_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1079_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1076_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1094_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1113_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1123_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1126_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1085_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1091_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1129_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1097_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1100_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1082_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1120_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1088_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1079_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1076_inst_req_1;
      WPIPE_Block2_start_1094_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1113_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1123_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1126_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1085_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1091_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1129_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1097_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1100_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1082_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1120_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1088_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1079_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1076_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add57_214 & conv322_1112 & add117_365 & add126_390 & add30_139 & add48_189 & add135_415 & add99_315 & add108_340 & add21_114 & conv324_1119 & add39_164 & add12_89 & add_64;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1135_inst WPIPE_Block3_start_1150_inst WPIPE_Block3_start_1147_inst WPIPE_Block3_start_1144_inst WPIPE_Block3_start_1132_inst WPIPE_Block3_start_1141_inst WPIPE_Block3_start_1138_inst WPIPE_Block3_start_1185_inst WPIPE_Block3_start_1156_inst WPIPE_Block3_start_1153_inst WPIPE_Block3_start_1182_inst WPIPE_Block3_start_1179_inst WPIPE_Block3_start_1176_inst WPIPE_Block3_start_1169_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1135_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1150_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1147_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1144_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1132_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1141_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1138_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1185_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1156_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1153_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1182_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1179_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1176_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1169_inst_req_0;
      WPIPE_Block3_start_1135_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1150_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1147_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1144_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1132_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1141_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1138_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1185_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1156_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1153_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1182_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1179_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1176_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1169_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1135_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1150_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1147_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1144_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1132_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1141_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1138_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1185_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1156_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1153_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1182_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1179_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1176_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1169_inst_req_1;
      WPIPE_Block3_start_1135_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1150_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1147_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1144_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1132_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1141_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1138_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1185_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1156_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1153_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1182_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1179_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1176_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1169_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add12_89 & add57_214 & add48_189 & add39_164 & add_64 & add30_139 & add21_114 & add135_415 & add108_340 & add99_315 & add126_390 & add117_365 & conv341_1175 & conv339_1168;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1309_inst WPIPE_ConvTranspose_output_pipe_1306_inst WPIPE_ConvTranspose_output_pipe_1303_inst WPIPE_ConvTranspose_output_pipe_1300_inst WPIPE_ConvTranspose_output_pipe_1297_inst WPIPE_ConvTranspose_output_pipe_1294_inst WPIPE_ConvTranspose_output_pipe_1291_inst WPIPE_ConvTranspose_output_pipe_1312_inst WPIPE_ConvTranspose_output_pipe_1453_inst WPIPE_ConvTranspose_output_pipe_1456_inst WPIPE_ConvTranspose_output_pipe_1459_inst WPIPE_ConvTranspose_output_pipe_1462_inst WPIPE_ConvTranspose_output_pipe_1465_inst WPIPE_ConvTranspose_output_pipe_1468_inst WPIPE_ConvTranspose_output_pipe_1471_inst WPIPE_ConvTranspose_output_pipe_1474_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1309_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1306_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1303_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1300_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1297_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1312_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1453_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1456_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1459_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1462_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1465_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1468_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1471_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1474_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1309_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1306_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1303_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1300_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1297_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1312_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1453_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1456_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1459_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1462_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1465_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1468_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1471_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1474_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1309_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1306_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1303_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1300_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1297_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1312_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1453_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1456_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1459_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1462_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1465_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1468_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1471_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1474_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1309_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1306_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1303_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1300_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1297_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1312_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1453_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1456_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1459_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1462_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1465_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1468_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1471_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1474_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv368_1230 & conv374_1240 & conv380_1250 & conv386_1260 & conv392_1270 & conv398_1280 & conv404_1290 & conv362_1220 & conv480_1452 & conv474_1442 & conv468_1432 & conv462_1422 & conv456_1412 & conv450_1402 & conv444_1392 & conv438_1382;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1214_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1214_inst_req_0;
      WPIPE_elapsed_time_pipe_1214_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1214_inst_req_1;
      WPIPE_elapsed_time_pipe_1214_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1213;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_968_call call_stmt_1203_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_968_call_req_0;
      reqL_unguarded(0) <= call_stmt_1203_call_req_0;
      call_stmt_968_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1203_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_968_call_req_1;
      reqR_unguarded(0) <= call_stmt_1203_call_req_1;
      call_stmt_968_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1203_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_968 <= data_out(127 downto 64);
      call354_1203 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3777_start: Boolean;
  signal convTransposeA_CP_3777_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1559_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1528_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1513_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1513_inst_ack_0 : boolean;
  signal type_cast_1548_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1559_inst_ack_0 : boolean;
  signal type_cast_1548_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1528_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1510_inst_ack_0 : boolean;
  signal type_cast_1548_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1544_inst_ack_0 : boolean;
  signal type_cast_1535_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1544_inst_req_0 : boolean;
  signal type_cast_1548_inst_ack_0 : boolean;
  signal type_cast_1535_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1528_inst_ack_1 : boolean;
  signal type_cast_1638_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1528_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1507_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1525_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1519_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1519_inst_ack_0 : boolean;
  signal phi_stmt_1820_req_1 : boolean;
  signal RPIPE_Block0_start_1525_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1510_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1513_inst_ack_1 : boolean;
  signal type_cast_1836_inst_ack_0 : boolean;
  signal type_cast_1826_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1525_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1513_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1510_inst_req_1 : boolean;
  signal type_cast_1836_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1544_inst_req_1 : boolean;
  signal type_cast_1617_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1544_inst_ack_1 : boolean;
  signal phi_stmt_1632_req_1 : boolean;
  signal type_cast_1826_inst_ack_1 : boolean;
  signal type_cast_1617_inst_ack_1 : boolean;
  signal type_cast_1638_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1516_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1507_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1516_inst_ack_0 : boolean;
  signal phi_stmt_1820_req_0 : boolean;
  signal type_cast_1836_inst_req_1 : boolean;
  signal type_cast_1638_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1525_inst_ack_1 : boolean;
  signal phi_stmt_1632_req_0 : boolean;
  signal RPIPE_Block0_start_1519_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1507_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1519_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1559_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1562_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1507_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1556_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1504_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1504_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1562_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1556_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1531_inst_req_0 : boolean;
  signal type_cast_1589_inst_req_0 : boolean;
  signal type_cast_1589_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1559_inst_ack_1 : boolean;
  signal phi_stmt_1618_req_0 : boolean;
  signal RPIPE_Block0_start_1522_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1531_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1562_inst_req_0 : boolean;
  signal type_cast_1535_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1516_inst_req_1 : boolean;
  signal type_cast_1535_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1562_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1522_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1556_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1504_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1516_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1531_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1504_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1556_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1510_inst_req_0 : boolean;
  signal type_cast_1836_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1531_inst_ack_1 : boolean;
  signal phi_stmt_1611_req_0 : boolean;
  signal phi_stmt_1611_req_1 : boolean;
  signal type_cast_1638_inst_ack_0 : boolean;
  signal type_cast_1838_inst_req_0 : boolean;
  signal type_cast_1838_inst_ack_0 : boolean;
  signal type_cast_1589_inst_req_1 : boolean;
  signal type_cast_1589_inst_ack_1 : boolean;
  signal type_cast_1593_inst_req_0 : boolean;
  signal type_cast_1593_inst_ack_0 : boolean;
  signal type_cast_1593_inst_req_1 : boolean;
  signal type_cast_1593_inst_ack_1 : boolean;
  signal phi_stmt_1827_req_1 : boolean;
  signal type_cast_1597_inst_req_0 : boolean;
  signal type_cast_1597_inst_ack_0 : boolean;
  signal type_cast_1832_inst_ack_1 : boolean;
  signal type_cast_1597_inst_req_1 : boolean;
  signal type_cast_1597_inst_ack_1 : boolean;
  signal phi_stmt_1827_req_0 : boolean;
  signal type_cast_1830_inst_ack_1 : boolean;
  signal type_cast_1830_inst_req_1 : boolean;
  signal type_cast_1832_inst_req_1 : boolean;
  signal type_cast_1601_inst_req_0 : boolean;
  signal type_cast_1601_inst_ack_0 : boolean;
  signal type_cast_1601_inst_req_1 : boolean;
  signal type_cast_1601_inst_ack_1 : boolean;
  signal type_cast_1826_inst_ack_0 : boolean;
  signal type_cast_1673_inst_req_0 : boolean;
  signal type_cast_1673_inst_ack_0 : boolean;
  signal type_cast_1832_inst_ack_0 : boolean;
  signal type_cast_1832_inst_req_0 : boolean;
  signal type_cast_1673_inst_req_1 : boolean;
  signal type_cast_1673_inst_ack_1 : boolean;
  signal type_cast_1830_inst_ack_0 : boolean;
  signal type_cast_1826_inst_req_0 : boolean;
  signal type_cast_1677_inst_req_0 : boolean;
  signal type_cast_1677_inst_ack_0 : boolean;
  signal type_cast_1677_inst_req_1 : boolean;
  signal type_cast_1677_inst_ack_1 : boolean;
  signal type_cast_1830_inst_req_0 : boolean;
  signal type_cast_1681_inst_req_0 : boolean;
  signal type_cast_1681_inst_ack_0 : boolean;
  signal type_cast_1681_inst_req_1 : boolean;
  signal type_cast_1681_inst_ack_1 : boolean;
  signal type_cast_1711_inst_req_0 : boolean;
  signal type_cast_1711_inst_ack_0 : boolean;
  signal type_cast_1711_inst_req_1 : boolean;
  signal type_cast_1711_inst_ack_1 : boolean;
  signal phi_stmt_1833_ack_0 : boolean;
  signal phi_stmt_1827_ack_0 : boolean;
  signal phi_stmt_1833_req_1 : boolean;
  signal type_cast_1838_inst_ack_1 : boolean;
  signal WPIPE_Block0_done_1849_inst_ack_0 : boolean;
  signal phi_stmt_1625_req_1 : boolean;
  signal type_cast_1838_inst_req_1 : boolean;
  signal type_cast_1631_inst_ack_1 : boolean;
  signal type_cast_1631_inst_req_1 : boolean;
  signal array_obj_ref_1717_index_offset_req_0 : boolean;
  signal array_obj_ref_1717_index_offset_ack_0 : boolean;
  signal array_obj_ref_1717_index_offset_req_1 : boolean;
  signal array_obj_ref_1717_index_offset_ack_1 : boolean;
  signal addr_of_1718_final_reg_req_0 : boolean;
  signal addr_of_1718_final_reg_ack_0 : boolean;
  signal WPIPE_Block0_done_1849_inst_ack_1 : boolean;
  signal addr_of_1718_final_reg_req_1 : boolean;
  signal addr_of_1718_final_reg_ack_1 : boolean;
  signal phi_stmt_1820_ack_0 : boolean;
  signal type_cast_1631_inst_ack_0 : boolean;
  signal type_cast_1631_inst_req_0 : boolean;
  signal phi_stmt_1632_ack_0 : boolean;
  signal phi_stmt_1625_req_0 : boolean;
  signal phi_stmt_1625_ack_0 : boolean;
  signal WPIPE_Block0_done_1849_inst_req_1 : boolean;
  signal phi_stmt_1618_ack_0 : boolean;
  signal type_cast_1617_inst_ack_0 : boolean;
  signal type_cast_1617_inst_req_0 : boolean;
  signal ptr_deref_1722_load_0_req_0 : boolean;
  signal ptr_deref_1722_load_0_ack_0 : boolean;
  signal ptr_deref_1722_load_0_req_1 : boolean;
  signal phi_stmt_1618_req_1 : boolean;
  signal ptr_deref_1722_load_0_ack_1 : boolean;
  signal phi_stmt_1833_req_0 : boolean;
  signal type_cast_1624_inst_ack_1 : boolean;
  signal phi_stmt_1611_ack_0 : boolean;
  signal type_cast_1624_inst_req_1 : boolean;
  signal type_cast_1624_inst_ack_0 : boolean;
  signal type_cast_1624_inst_req_0 : boolean;
  signal array_obj_ref_1740_index_offset_req_0 : boolean;
  signal array_obj_ref_1740_index_offset_ack_0 : boolean;
  signal array_obj_ref_1740_index_offset_req_1 : boolean;
  signal array_obj_ref_1740_index_offset_ack_1 : boolean;
  signal addr_of_1741_final_reg_req_0 : boolean;
  signal addr_of_1741_final_reg_ack_0 : boolean;
  signal addr_of_1741_final_reg_req_1 : boolean;
  signal addr_of_1741_final_reg_ack_1 : boolean;
  signal ptr_deref_1744_store_0_req_0 : boolean;
  signal ptr_deref_1744_store_0_ack_0 : boolean;
  signal ptr_deref_1744_store_0_req_1 : boolean;
  signal ptr_deref_1744_store_0_ack_1 : boolean;
  signal type_cast_1749_inst_req_0 : boolean;
  signal type_cast_1749_inst_ack_0 : boolean;
  signal type_cast_1749_inst_req_1 : boolean;
  signal type_cast_1749_inst_ack_1 : boolean;
  signal if_stmt_1762_branch_req_0 : boolean;
  signal if_stmt_1762_branch_ack_1 : boolean;
  signal if_stmt_1762_branch_ack_0 : boolean;
  signal type_cast_1790_inst_req_0 : boolean;
  signal type_cast_1790_inst_ack_0 : boolean;
  signal type_cast_1790_inst_req_1 : boolean;
  signal type_cast_1790_inst_ack_1 : boolean;
  signal type_cast_1806_inst_req_0 : boolean;
  signal type_cast_1806_inst_ack_0 : boolean;
  signal type_cast_1806_inst_req_1 : boolean;
  signal type_cast_1806_inst_ack_1 : boolean;
  signal if_stmt_1813_branch_req_0 : boolean;
  signal if_stmt_1813_branch_ack_1 : boolean;
  signal if_stmt_1813_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1849_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3777_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3777_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3777_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3777_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3777: Block -- control-path 
    signal convTransposeA_CP_3777_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3777_elements(0) <= convTransposeA_CP_3777_start;
    convTransposeA_CP_3777_symbol <= convTransposeA_CP_3777_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563__entry__
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/$entry
      -- CP-element group 0: 	 branch_block_stmt_1502/$entry
      -- CP-element group 0: 	 branch_block_stmt_1502/branch_block_stmt_1502__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Update/$entry
      -- 
    cr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(0), ack => type_cast_1548_inst_req_1); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(0), ack => type_cast_1535_inst_req_1); -- 
    rr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(0), ack => RPIPE_Block0_start_1504_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1502/merge_stmt_1819__exit__
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/assign_stmt_1845__entry__
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/assign_stmt_1845__exit__
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/assign_stmt_1845/$entry
      -- CP-element group 1: 	 branch_block_stmt_1502/assign_stmt_1845/$exit
      -- 
    cr_4585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1638_inst_req_1); -- 
    cr_4516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1617_inst_req_1); -- 
    rr_4580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1638_inst_req_0); -- 
    cr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1631_inst_req_1); -- 
    rr_4557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1631_inst_req_0); -- 
    rr_4511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1617_inst_req_0); -- 
    cr_4539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1624_inst_req_1); -- 
    rr_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(1), ack => type_cast_1624_inst_req_0); -- 
    convTransposeA_CP_3777_elements(1) <= convTransposeA_CP_3777_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Update/cr
      -- 
    ra_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1504_inst_ack_0, ack => convTransposeA_CP_3777_elements(2)); -- 
    cr_3830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(2), ack => RPIPE_Block0_start_1504_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1504_Update/ca
      -- 
    ca_3831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1504_inst_ack_1, ack => convTransposeA_CP_3777_elements(3)); -- 
    rr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(3), ack => RPIPE_Block0_start_1507_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Update/cr
      -- 
    ra_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1507_inst_ack_0, ack => convTransposeA_CP_3777_elements(4)); -- 
    cr_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(4), ack => RPIPE_Block0_start_1507_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1507_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Sample/rr
      -- 
    ca_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1507_inst_ack_1, ack => convTransposeA_CP_3777_elements(5)); -- 
    rr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(5), ack => RPIPE_Block0_start_1510_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Sample/$exit
      -- 
    ra_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1510_inst_ack_0, ack => convTransposeA_CP_3777_elements(6)); -- 
    cr_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(6), ack => RPIPE_Block0_start_1510_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1510_update_completed_
      -- 
    ca_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1510_inst_ack_1, ack => convTransposeA_CP_3777_elements(7)); -- 
    rr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(7), ack => RPIPE_Block0_start_1513_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Sample/$exit
      -- 
    ra_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1513_inst_ack_0, ack => convTransposeA_CP_3777_elements(8)); -- 
    cr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(8), ack => RPIPE_Block0_start_1513_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1513_update_completed_
      -- 
    ca_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1513_inst_ack_1, ack => convTransposeA_CP_3777_elements(9)); -- 
    rr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(9), ack => RPIPE_Block0_start_1516_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Update/cr
      -- 
    ra_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1516_inst_ack_0, ack => convTransposeA_CP_3777_elements(10)); -- 
    cr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(10), ack => RPIPE_Block0_start_1516_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1516_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_sample_start_
      -- 
    ca_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1516_inst_ack_1, ack => convTransposeA_CP_3777_elements(11)); -- 
    rr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(11), ack => RPIPE_Block0_start_1519_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Update/cr
      -- 
    ra_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1519_inst_ack_0, ack => convTransposeA_CP_3777_elements(12)); -- 
    cr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(12), ack => RPIPE_Block0_start_1519_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1519_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Sample/rr
      -- 
    ca_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1519_inst_ack_1, ack => convTransposeA_CP_3777_elements(13)); -- 
    rr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(13), ack => RPIPE_Block0_start_1522_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Update/cr
      -- 
    ra_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1522_inst_ack_0, ack => convTransposeA_CP_3777_elements(14)); -- 
    cr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(14), ack => RPIPE_Block0_start_1522_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1522_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Sample/$entry
      -- 
    ca_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1522_inst_ack_1, ack => convTransposeA_CP_3777_elements(15)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(15), ack => RPIPE_Block0_start_1525_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_update_start_
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1525_inst_ack_0, ack => convTransposeA_CP_3777_elements(16)); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(16), ack => RPIPE_Block0_start_1525_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1525_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Sample/$entry
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1525_inst_ack_1, ack => convTransposeA_CP_3777_elements(17)); -- 
    rr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(17), ack => RPIPE_Block0_start_1528_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Sample/$exit
      -- 
    ra_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1528_inst_ack_0, ack => convTransposeA_CP_3777_elements(18)); -- 
    cr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(18), ack => RPIPE_Block0_start_1528_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1528_update_completed_
      -- 
    ca_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1528_inst_ack_1, ack => convTransposeA_CP_3777_elements(19)); -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(19), ack => RPIPE_Block0_start_1531_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Update/cr
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1531_inst_ack_0, ack => convTransposeA_CP_3777_elements(20)); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(20), ack => RPIPE_Block0_start_1531_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1531_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_sample_start_
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1531_inst_ack_1, ack => convTransposeA_CP_3777_elements(21)); -- 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(21), ack => type_cast_1535_inst_req_0); -- 
    rr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(21), ack => RPIPE_Block0_start_1544_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_sample_completed_
      -- 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1535_inst_ack_0, ack => convTransposeA_CP_3777_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1535_Update/$exit
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1535_inst_ack_1, ack => convTransposeA_CP_3777_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Update/cr
      -- 
    ra_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1544_inst_ack_0, ack => convTransposeA_CP_3777_elements(24)); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(24), ack => RPIPE_Block0_start_1544_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1544_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Sample/rr
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1544_inst_ack_1, ack => convTransposeA_CP_3777_elements(25)); -- 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(25), ack => type_cast_1548_inst_req_0); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(25), ack => RPIPE_Block0_start_1556_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_sample_completed_
      -- 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1548_inst_ack_0, ack => convTransposeA_CP_3777_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/type_cast_1548_update_completed_
      -- 
    ca_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1548_inst_ack_1, ack => convTransposeA_CP_3777_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Update/cr
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1556_inst_ack_0, ack => convTransposeA_CP_3777_elements(28)); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(28), ack => RPIPE_Block0_start_1556_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1556_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_sample_start_
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1556_inst_ack_1, ack => convTransposeA_CP_3777_elements(29)); -- 
    rr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(29), ack => RPIPE_Block0_start_1559_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_update_start_
      -- 
    ra_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1559_inst_ack_0, ack => convTransposeA_CP_3777_elements(30)); -- 
    cr_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(30), ack => RPIPE_Block0_start_1559_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1559_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Sample/rr
      -- 
    ca_4027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1559_inst_ack_1, ack => convTransposeA_CP_3777_elements(31)); -- 
    rr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(31), ack => RPIPE_Block0_start_1562_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_update_start_
      -- 
    ra_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1562_inst_ack_0, ack => convTransposeA_CP_3777_elements(32)); -- 
    cr_4040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(32), ack => RPIPE_Block0_start_1562_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/RPIPE_Block0_start_1562_Update/ca
      -- 
    ca_4041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1562_inst_ack_1, ack => convTransposeA_CP_3777_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563/$exit
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608__entry__
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1505_to_assign_stmt_1563__exit__
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Update/cr
      -- 
    rr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1589_inst_req_0); -- 
    cr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1589_inst_req_1); -- 
    rr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1593_inst_req_0); -- 
    cr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1593_inst_req_1); -- 
    rr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1597_inst_req_0); -- 
    cr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1597_inst_req_1); -- 
    rr_4094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1601_inst_req_0); -- 
    cr_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(34), ack => type_cast_1601_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(23) & convTransposeA_CP_3777_elements(27) & convTransposeA_CP_3777_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Sample/$exit
      -- 
    ra_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_0, ack => convTransposeA_CP_3777_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1589_Update/ca
      -- 
    ca_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_1, ack => convTransposeA_CP_3777_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Sample/ra
      -- 
    ra_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1593_inst_ack_0, ack => convTransposeA_CP_3777_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1593_Update/ca
      -- 
    ca_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1593_inst_ack_1, ack => convTransposeA_CP_3777_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Sample/ra
      -- 
    ra_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_0, ack => convTransposeA_CP_3777_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1597_Update/ca
      -- 
    ca_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_1, ack => convTransposeA_CP_3777_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Sample/ra
      -- 
    ra_4095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_0, ack => convTransposeA_CP_3777_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/type_cast_1601_Update/ca
      -- 
    ca_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_1, ack => convTransposeA_CP_3777_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608__exit__
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1611/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1625/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1502/assign_stmt_1570_to_assign_stmt_1608/$exit
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1618/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1632/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(36) & convTransposeA_CP_3777_elements(38) & convTransposeA_CP_3777_elements(40) & convTransposeA_CP_3777_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Sample/ra
      -- 
    ra_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_0, ack => convTransposeA_CP_3777_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Update/ca
      -- 
    ca_4117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1673_inst_ack_1, ack => convTransposeA_CP_3777_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Sample/ra
      -- 
    ra_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1677_inst_ack_0, ack => convTransposeA_CP_3777_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Update/ca
      -- 
    ca_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1677_inst_ack_1, ack => convTransposeA_CP_3777_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Sample/ra
      -- 
    ra_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1681_inst_ack_0, ack => convTransposeA_CP_3777_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Update/ca
      -- 
    ca_4145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1681_inst_ack_1, ack => convTransposeA_CP_3777_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Sample/ra
      -- 
    ra_4154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_0, ack => convTransposeA_CP_3777_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Sample/req
      -- 
    ca_4159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_1, ack => convTransposeA_CP_3777_elements(51)); -- 
    req_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(51), ack => array_obj_ref_1717_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Sample/ack
      -- 
    ack_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1717_index_offset_ack_0, ack => convTransposeA_CP_3777_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_request/req
      -- 
    ack_4190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1717_index_offset_ack_1, ack => convTransposeA_CP_3777_elements(53)); -- 
    req_4199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(53), ack => addr_of_1718_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_request/ack
      -- 
    ack_4200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1718_final_reg_ack_0, ack => convTransposeA_CP_3777_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/word_access_start/word_0/rr
      -- 
    ack_4205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1718_final_reg_ack_1, ack => convTransposeA_CP_3777_elements(55)); -- 
    rr_4238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(55), ack => ptr_deref_1722_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Sample/word_access_start/word_0/ra
      -- 
    ra_4239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1722_load_0_ack_0, ack => convTransposeA_CP_3777_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/ptr_deref_1722_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/ptr_deref_1722_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/ptr_deref_1722_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/ptr_deref_1722_Merge/merge_ack
      -- 
    ca_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1722_load_0_ack_1, ack => convTransposeA_CP_3777_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Sample/req
      -- 
    req_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(58), ack => array_obj_ref_1740_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(45) & convTransposeA_CP_3777_elements(47) & convTransposeA_CP_3777_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Sample/ack
      -- 
    ack_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1740_index_offset_ack_0, ack => convTransposeA_CP_3777_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_request/req
      -- 
    ack_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1740_index_offset_ack_1, ack => convTransposeA_CP_3777_elements(60)); -- 
    req_4295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(60), ack => addr_of_1741_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_request/ack
      -- 
    ack_4296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1741_final_reg_ack_0, ack => convTransposeA_CP_3777_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_word_addrgen/root_register_ack
      -- 
    ack_4301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1741_final_reg_ack_1, ack => convTransposeA_CP_3777_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/ptr_deref_1744_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/ptr_deref_1744_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/ptr_deref_1744_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/ptr_deref_1744_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/word_access_start/word_0/rr
      -- 
    rr_4339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(63), ack => ptr_deref_1744_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(57) & convTransposeA_CP_3777_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Sample/word_access_start/word_0/ra
      -- 
    ra_4340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1744_store_0_ack_0, ack => convTransposeA_CP_3777_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/word_access_complete/word_0/ca
      -- 
    ca_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1744_store_0_ack_1, ack => convTransposeA_CP_3777_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Sample/ra
      -- 
    ra_4360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_0, ack => convTransposeA_CP_3777_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Update/ca
      -- 
    ca_4365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1749_inst_ack_1, ack => convTransposeA_CP_3777_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761__exit__
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762__entry__
      -- CP-element group 68: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/$exit
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1502/R_cmp_1763_place
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1502/if_stmt_1762_else_link/$entry
      -- 
    branch_req_4373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(68), ack => if_stmt_1762_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(52) & convTransposeA_CP_3777_elements(59) & convTransposeA_CP_3777_elements(65) & convTransposeA_CP_3777_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/merge_stmt_1768__exit__
      -- CP-element group 69: 	 branch_block_stmt_1502/assign_stmt_1774__entry__
      -- CP-element group 69: 	 branch_block_stmt_1502/assign_stmt_1774__exit__
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/merge_stmt_1768_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/merge_stmt_1768_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1502/merge_stmt_1768_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1502/merge_stmt_1768_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/if_stmt_1762_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1502/if_stmt_1762_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1502/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1502/assign_stmt_1774/$entry
      -- CP-element group 69: 	 branch_block_stmt_1502/assign_stmt_1774/$exit
      -- 
    if_choice_transition_4378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1762_branch_ack_1, ack => convTransposeA_CP_3777_elements(69)); -- 
    cr_4746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1826_inst_req_1); -- 
    rr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1836_inst_req_0); -- 
    cr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1836_inst_req_1); -- 
    cr_4723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1832_inst_req_1); -- 
    rr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1832_inst_req_0); -- 
    rr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(69), ack => type_cast_1826_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1502/merge_stmt_1776__exit__
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812__entry__
      -- CP-element group 70: 	 branch_block_stmt_1502/merge_stmt_1776_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1502/merge_stmt_1776_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1502/merge_stmt_1776_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1502/merge_stmt_1776_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1502/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/if_stmt_1762_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1502/if_stmt_1762_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1502/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Update/cr
      -- 
    else_choice_transition_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1762_branch_ack_0, ack => convTransposeA_CP_3777_elements(70)); -- 
    rr_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(70), ack => type_cast_1790_inst_req_0); -- 
    cr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(70), ack => type_cast_1790_inst_req_1); -- 
    cr_4417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(70), ack => type_cast_1806_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Sample/ra
      -- 
    ra_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1790_inst_ack_0, ack => convTransposeA_CP_3777_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1790_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Sample/rr
      -- 
    ca_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1790_inst_ack_1, ack => convTransposeA_CP_3777_elements(72)); -- 
    rr_4412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(72), ack => type_cast_1806_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Sample/ra
      -- 
    ra_4413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1806_inst_ack_0, ack => convTransposeA_CP_3777_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812__exit__
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813__entry__
      -- CP-element group 74: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/$exit
      -- CP-element group 74: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1502/assign_stmt_1782_to_assign_stmt_1812/type_cast_1806_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1502/R_cmp112_1814_place
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1502/if_stmt_1813_else_link/$entry
      -- 
    ca_4418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1806_inst_ack_1, ack => convTransposeA_CP_3777_elements(74)); -- 
    branch_req_4426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(74), ack => if_stmt_1813_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1502/assign_stmt_1852__entry__
      -- CP-element group 75: 	 branch_block_stmt_1502/merge_stmt_1847__exit__
      -- CP-element group 75: 	 branch_block_stmt_1502/merge_stmt_1847_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1502/merge_stmt_1847_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1502/merge_stmt_1847_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1502/merge_stmt_1847_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1502/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1502/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1502/if_stmt_1813_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1502/if_stmt_1813_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1502/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1502/assign_stmt_1852/$entry
      -- CP-element group 75: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Sample/req
      -- 
    if_choice_transition_4431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1813_branch_ack_1, ack => convTransposeA_CP_3777_elements(75)); -- 
    req_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(75), ack => WPIPE_Block0_done_1849_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1820/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1502/if_stmt_1813_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1502/if_stmt_1813_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123
      -- 
    else_choice_transition_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1813_branch_ack_0, ack => convTransposeA_CP_3777_elements(76)); -- 
    rr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1838_inst_req_0); -- 
    cr_4666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1830_inst_req_1); -- 
    rr_4661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1830_inst_req_0); -- 
    cr_4643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(76), ack => type_cast_1838_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Sample/$exit
      -- 
    ack_4452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1849_inst_ack_0, ack => convTransposeA_CP_3777_elements(77)); -- 
    req_4456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(77), ack => WPIPE_Block0_done_1849_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1502/merge_stmt_1854__exit__
      -- CP-element group 78: 	 branch_block_stmt_1502/assign_stmt_1852__exit__
      -- CP-element group 78: 	 branch_block_stmt_1502/return__
      -- CP-element group 78: 	 branch_block_stmt_1502/branch_block_stmt_1502__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1502/$exit
      -- CP-element group 78: 	 branch_block_stmt_1502/merge_stmt_1854_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1502/merge_stmt_1854_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1502/merge_stmt_1854_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1502/merge_stmt_1854_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1502/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1502/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1502/assign_stmt_1852/$exit
      -- CP-element group 78: 	 branch_block_stmt_1502/assign_stmt_1852/WPIPE_Block0_done_1849_update_completed_
      -- 
    ack_4457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1849_inst_ack_1, ack => convTransposeA_CP_3777_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1611/$exit
      -- CP-element group 79: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1615_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_req
      -- 
    phi_stmt_1611_req_4468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1611_req_4468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(79), ack => phi_stmt_1611_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1618/$exit
      -- CP-element group 80: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_req
      -- CP-element group 80: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1622_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$exit
      -- 
    phi_stmt_1618_req_4476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1618_req_4476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(80), ack => phi_stmt_1618_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1625/$exit
      -- CP-element group 81: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_req
      -- CP-element group 81: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1629_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/$exit
      -- 
    phi_stmt_1625_req_4484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1625_req_4484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(81), ack => phi_stmt_1625_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1636_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_req
      -- CP-element group 82: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/phi_stmt_1632/$exit
      -- 
    phi_stmt_1632_req_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1632_req_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(82), ack => phi_stmt_1632_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(43), ack => convTransposeA_CP_3777_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1502/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(79) & convTransposeA_CP_3777_elements(80) & convTransposeA_CP_3777_elements(81) & convTransposeA_CP_3777_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Sample/$exit
      -- 
    ra_4512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_0, ack => convTransposeA_CP_3777_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Update/ca
      -- CP-element group 85: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/Update/$exit
      -- 
    ca_4517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_1, ack => convTransposeA_CP_3777_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/$exit
      -- CP-element group 86: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_req
      -- CP-element group 86: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/$exit
      -- CP-element group 86: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1611/phi_stmt_1611_sources/type_cast_1617/SplitProtocol/$exit
      -- 
    phi_stmt_1611_req_4518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1611_req_4518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(86), ack => phi_stmt_1611_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(84) & convTransposeA_CP_3777_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Sample/$exit
      -- 
    ra_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1624_inst_ack_0, ack => convTransposeA_CP_3777_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Update/ca
      -- CP-element group 88: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/Update/$exit
      -- 
    ca_4540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1624_inst_ack_1, ack => convTransposeA_CP_3777_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_req
      -- CP-element group 89: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/type_cast_1624/$exit
      -- CP-element group 89: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/phi_stmt_1618_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1618/$exit
      -- 
    phi_stmt_1618_req_4541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1618_req_4541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(89), ack => phi_stmt_1618_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(87) & convTransposeA_CP_3777_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Sample/$exit
      -- 
    ra_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1631_inst_ack_0, ack => convTransposeA_CP_3777_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/Update/$exit
      -- 
    ca_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1631_inst_ack_1, ack => convTransposeA_CP_3777_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_req
      -- CP-element group 92: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1631/$exit
      -- CP-element group 92: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1625/$exit
      -- 
    phi_stmt_1625_req_4564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1625_req_4564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(92), ack => phi_stmt_1625_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(90) & convTransposeA_CP_3777_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/ra
      -- 
    ra_4581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_0, ack => convTransposeA_CP_3777_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/$exit
      -- 
    ca_4586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_1, ack => convTransposeA_CP_3777_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_req
      -- CP-element group 95: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/$exit
      -- CP-element group 95: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1632/$exit
      -- 
    phi_stmt_1632_req_4587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1632_req_4587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(95), ack => phi_stmt_1632_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(93) & convTransposeA_CP_3777_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1502/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(86) & convTransposeA_CP_3777_elements(89) & convTransposeA_CP_3777_elements(92) & convTransposeA_CP_3777_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1502/merge_stmt_1610_PhiAck/$entry
      -- CP-element group 97: 	 branch_block_stmt_1502/merge_stmt_1610_PhiReqMerge
      -- 
    convTransposeA_CP_3777_elements(97) <= OrReduce(convTransposeA_CP_3777_elements(83) & convTransposeA_CP_3777_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1502/merge_stmt_1610_PhiAck/phi_stmt_1611_ack
      -- 
    phi_stmt_1611_ack_4592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1611_ack_0, ack => convTransposeA_CP_3777_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1502/merge_stmt_1610_PhiAck/phi_stmt_1618_ack
      -- 
    phi_stmt_1618_ack_4593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1618_ack_0, ack => convTransposeA_CP_3777_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1502/merge_stmt_1610_PhiAck/phi_stmt_1625_ack
      -- 
    phi_stmt_1625_ack_4594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1625_ack_0, ack => convTransposeA_CP_3777_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1502/merge_stmt_1610_PhiAck/phi_stmt_1632_ack
      -- 
    phi_stmt_1632_ack_4595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1632_ack_0, ack => convTransposeA_CP_3777_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1502/merge_stmt_1610__exit__
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761__entry__
      -- CP-element group 102: 	 branch_block_stmt_1502/merge_stmt_1610_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1673_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1677_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1681_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1711_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1717_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1718_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1722_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/array_obj_ref_1740_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/addr_of_1741_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/ptr_deref_1744_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1502/assign_stmt_1645_to_assign_stmt_1761/type_cast_1749_Update/cr
      -- 
    rr_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1673_inst_req_0); -- 
    cr_4116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1673_inst_req_1); -- 
    rr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1677_inst_req_0); -- 
    cr_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1677_inst_req_1); -- 
    rr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1681_inst_req_0); -- 
    cr_4144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1681_inst_req_1); -- 
    rr_4153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1711_inst_req_0); -- 
    cr_4158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1711_inst_req_1); -- 
    req_4189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => array_obj_ref_1717_index_offset_req_1); -- 
    req_4204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => addr_of_1718_final_reg_req_1); -- 
    cr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => ptr_deref_1722_load_0_req_1); -- 
    req_4285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => array_obj_ref_1740_index_offset_req_1); -- 
    req_4300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => addr_of_1741_final_reg_req_1); -- 
    cr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => ptr_deref_1744_store_0_req_1); -- 
    rr_4359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1749_inst_req_0); -- 
    cr_4364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(102), ack => type_cast_1749_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(98) & convTransposeA_CP_3777_elements(99) & convTransposeA_CP_3777_elements(100) & convTransposeA_CP_3777_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Sample/ra
      -- 
    ra_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1838_inst_ack_0, ack => convTransposeA_CP_3777_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/Update/$exit
      -- 
    ca_4644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1838_inst_ack_1, ack => convTransposeA_CP_3777_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1838/$exit
      -- CP-element group 105: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/$exit
      -- CP-element group 105: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_req
      -- 
    phi_stmt_1833_req_4645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1833_req_4645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(105), ack => phi_stmt_1833_req_1); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(103) & convTransposeA_CP_3777_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Sample/$exit
      -- 
    ra_4662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_0, ack => convTransposeA_CP_3777_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/ca
      -- CP-element group 107: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/Update/$exit
      -- 
    ca_4667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_1, ack => convTransposeA_CP_3777_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_req
      -- CP-element group 108: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1830/$exit
      -- CP-element group 108: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1827/$exit
      -- 
    phi_stmt_1827_req_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1827_req_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(108), ack => phi_stmt_1827_req_0); -- 
    convTransposeA_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(106) & convTransposeA_CP_3777_elements(107);
      gj_convTransposeA_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  output  delay-element  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_req
      -- CP-element group 109: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1824_konst_delay_trans
      -- CP-element group 109: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1820/$exit
      -- 
    phi_stmt_1820_req_4676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1820_req_4676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(109), ack => phi_stmt_1820_req_0); -- 
    -- Element group convTransposeA_CP_3777_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => convTransposeA_CP_3777_elements(76), ack => convTransposeA_CP_3777_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1502/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(105) & convTransposeA_CP_3777_elements(108) & convTransposeA_CP_3777_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Sample/ra
      -- 
    ra_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1836_inst_ack_0, ack => convTransposeA_CP_3777_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/Update/$exit
      -- 
    ca_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1836_inst_ack_1, ack => convTransposeA_CP_3777_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/$exit
      -- CP-element group 113: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1836/$exit
      -- CP-element group 113: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_req
      -- CP-element group 113: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$exit
      -- 
    phi_stmt_1833_req_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1833_req_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(113), ack => phi_stmt_1833_req_0); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(111) & convTransposeA_CP_3777_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Sample/$exit
      -- 
    ra_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_0, ack => convTransposeA_CP_3777_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/Update/$exit
      -- 
    ca_4724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_1, ack => convTransposeA_CP_3777_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_req
      -- CP-element group 116: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/type_cast_1832/$exit
      -- CP-element group 116: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/phi_stmt_1827_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1827/$exit
      -- 
    phi_stmt_1827_req_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1827_req_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(116), ack => phi_stmt_1827_req_1); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(114) & convTransposeA_CP_3777_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Sample/$exit
      -- 
    ra_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_0, ack => convTransposeA_CP_3777_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Update/ca
      -- CP-element group 118: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/Update/$exit
      -- 
    ca_4747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_1, ack => convTransposeA_CP_3777_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_req
      -- CP-element group 119: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/$exit
      -- CP-element group 119: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/$exit
      -- CP-element group 119: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1820/phi_stmt_1820_sources/type_cast_1826/SplitProtocol/$exit
      -- 
    phi_stmt_1820_req_4748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1820_req_4748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3777_elements(119), ack => phi_stmt_1820_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(117) & convTransposeA_CP_3777_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1502/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(113) & convTransposeA_CP_3777_elements(116) & convTransposeA_CP_3777_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1502/merge_stmt_1819_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_1502/merge_stmt_1819_PhiReqMerge
      -- 
    convTransposeA_CP_3777_elements(121) <= OrReduce(convTransposeA_CP_3777_elements(110) & convTransposeA_CP_3777_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1502/merge_stmt_1819_PhiAck/phi_stmt_1820_ack
      -- 
    phi_stmt_1820_ack_4753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1820_ack_0, ack => convTransposeA_CP_3777_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1502/merge_stmt_1819_PhiAck/phi_stmt_1827_ack
      -- 
    phi_stmt_1827_ack_4754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1827_ack_0, ack => convTransposeA_CP_3777_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1502/merge_stmt_1819_PhiAck/phi_stmt_1833_ack
      -- 
    phi_stmt_1833_ack_4755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1833_ack_0, ack => convTransposeA_CP_3777_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1502/merge_stmt_1819_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3777_elements(122) & convTransposeA_CP_3777_elements(123) & convTransposeA_CP_3777_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3777_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1739_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1739_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1716_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1716_scaled : std_logic_vector(13 downto 0);
    signal add41_1570 : std_logic_vector(15 downto 0);
    signal add54_1581 : std_logic_vector(15 downto 0);
    signal add73_1692 : std_logic_vector(63 downto 0);
    signal add75_1702 : std_logic_vector(63 downto 0);
    signal add86_1756 : std_logic_vector(31 downto 0);
    signal add93_1774 : std_logic_vector(15 downto 0);
    signal add_1554 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1650 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1717_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1740_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1740_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1740_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1740_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1740_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1740_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1719 : std_logic_vector(31 downto 0);
    signal arrayidx82_1742 : std_logic_vector(31 downto 0);
    signal call11_1523 : std_logic_vector(15 downto 0);
    signal call13_1526 : std_logic_vector(15 downto 0);
    signal call14_1529 : std_logic_vector(15 downto 0);
    signal call15_1532 : std_logic_vector(15 downto 0);
    signal call16_1545 : std_logic_vector(15 downto 0);
    signal call18_1557 : std_logic_vector(15 downto 0);
    signal call1_1508 : std_logic_vector(15 downto 0);
    signal call20_1560 : std_logic_vector(15 downto 0);
    signal call22_1563 : std_logic_vector(15 downto 0);
    signal call3_1511 : std_logic_vector(15 downto 0);
    signal call5_1514 : std_logic_vector(15 downto 0);
    signal call7_1517 : std_logic_vector(15 downto 0);
    signal call9_1520 : std_logic_vector(15 downto 0);
    signal call_1505 : std_logic_vector(15 downto 0);
    signal cmp101_1787 : std_logic_vector(0 downto 0);
    signal cmp112_1812 : std_logic_vector(0 downto 0);
    signal cmp_1761 : std_logic_vector(0 downto 0);
    signal conv107_1807 : std_logic_vector(31 downto 0);
    signal conv110_1602 : std_logic_vector(31 downto 0);
    signal conv17_1549 : std_logic_vector(31 downto 0);
    signal conv61_1674 : std_logic_vector(63 downto 0);
    signal conv64_1590 : std_logic_vector(63 downto 0);
    signal conv66_1678 : std_logic_vector(63 downto 0);
    signal conv69_1594 : std_logic_vector(63 downto 0);
    signal conv71_1682 : std_logic_vector(63 downto 0);
    signal conv85_1750 : std_logic_vector(31 downto 0);
    signal conv89_1598 : std_logic_vector(31 downto 0);
    signal conv_1536 : std_logic_vector(31 downto 0);
    signal idxprom81_1735 : std_logic_vector(63 downto 0);
    signal idxprom_1712 : std_logic_vector(63 downto 0);
    signal inc105_1791 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1796 : std_logic_vector(15 downto 0);
    signal inc_1782 : std_logic_vector(15 downto 0);
    signal indvar_1611 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1845 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1833 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1632 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1827 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1625 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1803 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1820 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1618 : std_logic_vector(15 downto 0);
    signal mul50_1665 : std_logic_vector(15 downto 0);
    signal mul72_1687 : std_logic_vector(63 downto 0);
    signal mul74_1697 : std_logic_vector(63 downto 0);
    signal mul_1655 : std_logic_vector(15 downto 0);
    signal ptr_deref_1722_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1722_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1722_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1722_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1722_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1744_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1744_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1744_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1744_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1744_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1744_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1542 : std_logic_vector(31 downto 0);
    signal shr111126_1608 : std_logic_vector(31 downto 0);
    signal shr80_1729 : std_logic_vector(63 downto 0);
    signal shr_1708 : std_logic_vector(31 downto 0);
    signal sub44_1660 : std_logic_vector(15 downto 0);
    signal sub57_1586 : std_logic_vector(15 downto 0);
    signal sub58_1670 : std_logic_vector(15 downto 0);
    signal sub_1575 : std_logic_vector(15 downto 0);
    signal tmp1_1645 : std_logic_vector(31 downto 0);
    signal tmp78_1723 : std_logic_vector(63 downto 0);
    signal type_cast_1540_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1568_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1579_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1606_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1615_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1617_wire : std_logic_vector(31 downto 0);
    signal type_cast_1622_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1624_wire : std_logic_vector(15 downto 0);
    signal type_cast_1629_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1631_wire : std_logic_vector(15 downto 0);
    signal type_cast_1636_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1638_wire : std_logic_vector(15 downto 0);
    signal type_cast_1643_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1706_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1727_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1733_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1772_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1780_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1800_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1824_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1826_wire : std_logic_vector(15 downto 0);
    signal type_cast_1830_wire : std_logic_vector(15 downto 0);
    signal type_cast_1832_wire : std_logic_vector(15 downto 0);
    signal type_cast_1836_wire : std_logic_vector(15 downto 0);
    signal type_cast_1838_wire : std_logic_vector(15 downto 0);
    signal type_cast_1843_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1851_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1717_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1717_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1717_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1717_resized_base_address <= "00000000000000";
    array_obj_ref_1740_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1740_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1740_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1740_resized_base_address <= "00000000000000";
    ptr_deref_1722_word_offset_0 <= "00000000000000";
    ptr_deref_1744_word_offset_0 <= "00000000000000";
    type_cast_1540_wire_constant <= "00000000000000000000000000010000";
    type_cast_1568_wire_constant <= "1111111111111111";
    type_cast_1579_wire_constant <= "1111111111111111";
    type_cast_1606_wire_constant <= "00000000000000000000000000000010";
    type_cast_1615_wire_constant <= "00000000000000000000000000000000";
    type_cast_1622_wire_constant <= "0000000000000000";
    type_cast_1629_wire_constant <= "0000000000000000";
    type_cast_1636_wire_constant <= "0000000000000000";
    type_cast_1643_wire_constant <= "00000000000000000000000000000100";
    type_cast_1706_wire_constant <= "00000000000000000000000000000010";
    type_cast_1727_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1733_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1754_wire_constant <= "00000000000000000000000000000100";
    type_cast_1772_wire_constant <= "0000000000000100";
    type_cast_1780_wire_constant <= "0000000000000001";
    type_cast_1800_wire_constant <= "0000000000000000";
    type_cast_1824_wire_constant <= "0000000000000000";
    type_cast_1843_wire_constant <= "00000000000000000000000000000001";
    type_cast_1851_wire_constant <= "0000000000000001";
    phi_stmt_1611: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1615_wire_constant & type_cast_1617_wire;
      req <= phi_stmt_1611_req_0 & phi_stmt_1611_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1611",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1611_ack_0,
          idata => idata,
          odata => indvar_1611,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1611
    phi_stmt_1618: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1622_wire_constant & type_cast_1624_wire;
      req <= phi_stmt_1618_req_0 & phi_stmt_1618_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1618",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1618_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1618,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1618
    phi_stmt_1625: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1629_wire_constant & type_cast_1631_wire;
      req <= phi_stmt_1625_req_0 & phi_stmt_1625_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1625",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1625_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1625,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1625
    phi_stmt_1632: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1636_wire_constant & type_cast_1638_wire;
      req <= phi_stmt_1632_req_0 & phi_stmt_1632_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1632",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1632_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1632,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1632
    phi_stmt_1820: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1824_wire_constant & type_cast_1826_wire;
      req <= phi_stmt_1820_req_0 & phi_stmt_1820_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1820",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1820_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1820,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1820
    phi_stmt_1827: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1830_wire & type_cast_1832_wire;
      req <= phi_stmt_1827_req_0 & phi_stmt_1827_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1827",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1827_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1827
    phi_stmt_1833: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1836_wire & type_cast_1838_wire;
      req <= phi_stmt_1833_req_0 & phi_stmt_1833_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1833",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1833_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1833,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1833
    -- flow-through select operator MUX_1802_inst
    input_dim1x_x2_1803 <= type_cast_1800_wire_constant when (cmp101_1787(0) /=  '0') else inc_1782;
    addr_of_1718_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1718_final_reg_req_0;
      addr_of_1718_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1718_final_reg_req_1;
      addr_of_1718_final_reg_ack_1<= rack(0);
      addr_of_1718_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1718_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1717_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1741_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1741_final_reg_req_0;
      addr_of_1741_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1741_final_reg_req_1;
      addr_of_1741_final_reg_ack_1<= rack(0);
      addr_of_1741_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1741_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1740_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1535_inst_req_0;
      type_cast_1535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1535_inst_req_1;
      type_cast_1535_inst_ack_1<= rack(0);
      type_cast_1535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1532,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1548_inst_req_0;
      type_cast_1548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1548_inst_req_1;
      type_cast_1548_inst_ack_1<= rack(0);
      type_cast_1548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1589_inst_req_0;
      type_cast_1589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1589_inst_req_1;
      type_cast_1589_inst_ack_1<= rack(0);
      type_cast_1589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1563,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1593_inst_req_0;
      type_cast_1593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1593_inst_req_1;
      type_cast_1593_inst_ack_1<= rack(0);
      type_cast_1593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1560,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1597_inst_req_0;
      type_cast_1597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1597_inst_req_1;
      type_cast_1597_inst_ack_1<= rack(0);
      type_cast_1597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1601_inst_req_0;
      type_cast_1601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1601_inst_req_1;
      type_cast_1601_inst_ack_1<= rack(0);
      type_cast_1601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1617_inst_req_0;
      type_cast_1617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1617_inst_req_1;
      type_cast_1617_inst_ack_1<= rack(0);
      type_cast_1617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1845,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1617_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1624_inst_req_0;
      type_cast_1624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1624_inst_req_1;
      type_cast_1624_inst_ack_1<= rack(0);
      type_cast_1624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1624_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1631_inst_req_0;
      type_cast_1631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1631_inst_req_1;
      type_cast_1631_inst_ack_1<= rack(0);
      type_cast_1631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1827,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1631_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1638_inst_req_0;
      type_cast_1638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1638_inst_req_1;
      type_cast_1638_inst_ack_1<= rack(0);
      type_cast_1638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1638_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1673_inst_req_0;
      type_cast_1673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1673_inst_req_1;
      type_cast_1673_inst_ack_1<= rack(0);
      type_cast_1673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1677_inst_req_0;
      type_cast_1677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1677_inst_req_1;
      type_cast_1677_inst_ack_1<= rack(0);
      type_cast_1677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1681_inst_req_0;
      type_cast_1681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1681_inst_req_1;
      type_cast_1681_inst_ack_1<= rack(0);
      type_cast_1681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1711_inst_req_0;
      type_cast_1711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1711_inst_req_1;
      type_cast_1711_inst_ack_1<= rack(0);
      type_cast_1711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1712,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1749_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1749_inst_req_0;
      type_cast_1749_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1749_inst_req_1;
      type_cast_1749_inst_ack_1<= rack(0);
      type_cast_1749_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1749_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1750,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1790_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1790_inst_req_0;
      type_cast_1790_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1790_inst_req_1;
      type_cast_1790_inst_ack_1<= rack(0);
      type_cast_1790_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1790_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1787,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1791,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1806_inst_req_0;
      type_cast_1806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1806_inst_req_1;
      type_cast_1806_inst_ack_1<= rack(0);
      type_cast_1806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1826_inst_req_0;
      type_cast_1826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1826_inst_req_1;
      type_cast_1826_inst_ack_1<= rack(0);
      type_cast_1826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1774,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1826_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1830_inst_req_0;
      type_cast_1830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1830_inst_req_1;
      type_cast_1830_inst_ack_1<= rack(0);
      type_cast_1830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1830_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1832_inst_req_0;
      type_cast_1832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1832_inst_req_1;
      type_cast_1832_inst_ack_1<= rack(0);
      type_cast_1832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1832_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1836_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1836_inst_req_0;
      type_cast_1836_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1836_inst_req_1;
      type_cast_1836_inst_ack_1<= rack(0);
      type_cast_1836_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1836_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1836_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1838_inst_req_0;
      type_cast_1838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1838_inst_req_1;
      type_cast_1838_inst_ack_1<= rack(0);
      type_cast_1838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1838_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1717_index_1_rename
    process(R_idxprom_1716_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1716_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1716_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1717_index_1_resize
    process(idxprom_1712) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1712;
      ov := iv(13 downto 0);
      R_idxprom_1716_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1717_root_address_inst
    process(array_obj_ref_1717_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1717_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1717_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1740_index_1_rename
    process(R_idxprom81_1739_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1739_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1739_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1740_index_1_resize
    process(idxprom81_1735) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1735;
      ov := iv(13 downto 0);
      R_idxprom81_1739_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1740_root_address_inst
    process(array_obj_ref_1740_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1740_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1740_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1722_addr_0
    process(ptr_deref_1722_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1722_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1722_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1722_base_resize
    process(arrayidx77_1719) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1719;
      ov := iv(13 downto 0);
      ptr_deref_1722_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1722_gather_scatter
    process(ptr_deref_1722_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1722_data_0;
      ov(63 downto 0) := iv;
      tmp78_1723 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1722_root_address_inst
    process(ptr_deref_1722_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1722_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1722_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_addr_0
    process(ptr_deref_1744_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1744_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1744_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_base_resize
    process(arrayidx82_1742) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1742;
      ov := iv(13 downto 0);
      ptr_deref_1744_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_gather_scatter
    process(tmp78_1723) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1723;
      ov(63 downto 0) := iv;
      ptr_deref_1744_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_root_address_inst
    process(ptr_deref_1744_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1744_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1744_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1762_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1761;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1762_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1762_branch_req_0,
          ack0 => if_stmt_1762_branch_ack_0,
          ack1 => if_stmt_1762_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1813_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1812;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1813_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1813_branch_req_0,
          ack0 => if_stmt_1813_branch_ack_0,
          ack1 => if_stmt_1813_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1569_inst
    process(call7_1517) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1517, type_cast_1568_wire_constant, tmp_var);
      add41_1570 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1580_inst
    process(call9_1520) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1520, type_cast_1579_wire_constant, tmp_var);
      add54_1581 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1659_inst
    process(sub_1575, mul_1655) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1575, mul_1655, tmp_var);
      sub44_1660 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1669_inst
    process(sub57_1586, mul50_1665) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1586, mul50_1665, tmp_var);
      sub58_1670 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1773_inst
    process(input_dim2x_x1_1618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1618, type_cast_1772_wire_constant, tmp_var);
      add93_1774 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1781_inst
    process(input_dim1x_x1_1625) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1625, type_cast_1780_wire_constant, tmp_var);
      inc_1782 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1795_inst
    process(inc105_1791, input_dim0x_x2_1632) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1791, input_dim0x_x2_1632, tmp_var);
      inc105x_xinput_dim0x_x2_1796 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1649_inst
    process(add_1554, tmp1_1645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1554, tmp1_1645, tmp_var);
      add_src_0x_x0_1650 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1755_inst
    process(conv85_1750) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1750, type_cast_1754_wire_constant, tmp_var);
      add86_1756 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1844_inst
    process(indvar_1611) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1611, type_cast_1843_wire_constant, tmp_var);
      indvarx_xnext_1845 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1691_inst
    process(mul72_1687, conv66_1678) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1687, conv66_1678, tmp_var);
      add73_1692 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1701_inst
    process(mul74_1697, conv61_1674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1697, conv61_1674, tmp_var);
      add75_1702 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1734_inst
    process(shr80_1729) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1729, type_cast_1733_wire_constant, tmp_var);
      idxprom81_1735 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1786_inst
    process(inc_1782, call1_1508) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1782, call1_1508, tmp_var);
      cmp101_1787 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1811_inst
    process(conv107_1807, shr111126_1608) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1807, shr111126_1608, tmp_var);
      cmp112_1812 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1607_inst
    process(conv110_1602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1602, type_cast_1606_wire_constant, tmp_var);
      shr111126_1608 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1707_inst
    process(add_src_0x_x0_1650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1650, type_cast_1706_wire_constant, tmp_var);
      shr_1708 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1728_inst
    process(add75_1702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1702, type_cast_1727_wire_constant, tmp_var);
      shr80_1729 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1654_inst
    process(input_dim0x_x2_1632, call13_1526) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1632, call13_1526, tmp_var);
      mul_1655 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1664_inst
    process(input_dim1x_x1_1625, call13_1526) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1625, call13_1526, tmp_var);
      mul50_1665 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1644_inst
    process(indvar_1611) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1611, type_cast_1643_wire_constant, tmp_var);
      tmp1_1645 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1686_inst
    process(conv71_1682, conv69_1594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1682, conv69_1594, tmp_var);
      mul72_1687 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1696_inst
    process(add73_1692, conv64_1590) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1692, conv64_1590, tmp_var);
      mul74_1697 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1553_inst
    process(shl_1542, conv17_1549) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1542, conv17_1549, tmp_var);
      add_1554 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1541_inst
    process(conv_1536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1536, type_cast_1540_wire_constant, tmp_var);
      shl_1542 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1574_inst
    process(add41_1570, call14_1529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1570, call14_1529, tmp_var);
      sub_1575 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1585_inst
    process(add54_1581, call14_1529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1581, call14_1529, tmp_var);
      sub57_1586 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1760_inst
    process(add86_1756, conv89_1598) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1756, conv89_1598, tmp_var);
      cmp_1761 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1717_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1716_scaled;
      array_obj_ref_1717_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1717_index_offset_req_0;
      array_obj_ref_1717_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1717_index_offset_req_1;
      array_obj_ref_1717_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1740_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1739_scaled;
      array_obj_ref_1740_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1740_index_offset_req_0;
      array_obj_ref_1740_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1740_index_offset_req_1;
      array_obj_ref_1740_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1722_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1722_load_0_req_0;
      ptr_deref_1722_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1722_load_0_req_1;
      ptr_deref_1722_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1722_word_address_0;
      ptr_deref_1722_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1744_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1744_store_0_req_0;
      ptr_deref_1744_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1744_store_0_req_1;
      ptr_deref_1744_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1744_word_address_0;
      data_in <= ptr_deref_1744_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1510_inst RPIPE_Block0_start_1507_inst RPIPE_Block0_start_1513_inst RPIPE_Block0_start_1528_inst RPIPE_Block0_start_1504_inst RPIPE_Block0_start_1556_inst RPIPE_Block0_start_1516_inst RPIPE_Block0_start_1519_inst RPIPE_Block0_start_1531_inst RPIPE_Block0_start_1559_inst RPIPE_Block0_start_1522_inst RPIPE_Block0_start_1544_inst RPIPE_Block0_start_1562_inst RPIPE_Block0_start_1525_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1510_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1507_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1513_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1528_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1504_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1556_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1516_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1519_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1531_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1559_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1522_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1544_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1562_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1525_inst_req_0;
      RPIPE_Block0_start_1510_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1507_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1513_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1528_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1504_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1556_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1516_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1519_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1531_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1559_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1522_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1544_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1562_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1525_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1510_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1507_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1513_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1528_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1504_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1556_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1516_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1519_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1531_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1559_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1522_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1544_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1562_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1525_inst_req_1;
      RPIPE_Block0_start_1510_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1507_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1513_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1528_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1504_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1556_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1516_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1519_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1531_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1559_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1522_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1544_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1562_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1525_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call3_1511 <= data_out(223 downto 208);
      call1_1508 <= data_out(207 downto 192);
      call5_1514 <= data_out(191 downto 176);
      call14_1529 <= data_out(175 downto 160);
      call_1505 <= data_out(159 downto 144);
      call18_1557 <= data_out(143 downto 128);
      call7_1517 <= data_out(127 downto 112);
      call9_1520 <= data_out(111 downto 96);
      call15_1532 <= data_out(95 downto 80);
      call20_1560 <= data_out(79 downto 64);
      call11_1523 <= data_out(63 downto 48);
      call16_1545 <= data_out(47 downto 32);
      call22_1563 <= data_out(31 downto 16);
      call13_1526 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1849_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1849_inst_req_0;
      WPIPE_Block0_done_1849_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1849_inst_req_1;
      WPIPE_Block0_done_1849_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1851_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4772_start: Boolean;
  signal convTransposeB_CP_4772_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1878_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1900_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1881_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1881_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1878_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1863_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1875_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1878_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1881_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1869_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1869_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1860_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1860_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1872_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1866_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1860_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1866_inst_ack_0 : boolean;
  signal type_cast_2187_inst_req_1 : boolean;
  signal type_cast_2187_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1900_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1912_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1912_inst_ack_1 : boolean;
  signal type_cast_1904_inst_ack_0 : boolean;
  signal type_cast_1904_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1912_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1884_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1884_inst_req_1 : boolean;
  signal type_cast_1951_inst_ack_0 : boolean;
  signal type_cast_2187_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1878_inst_req_1 : boolean;
  signal phi_stmt_1973_ack_0 : boolean;
  signal RPIPE_Block1_start_1918_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1918_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1875_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1915_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1915_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1900_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1863_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1875_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1912_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1915_inst_ack_1 : boolean;
  signal phi_stmt_2181_req_1 : boolean;
  signal RPIPE_Block1_start_1884_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1875_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1869_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1884_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1881_inst_ack_0 : boolean;
  signal type_cast_1951_inst_req_0 : boolean;
  signal type_cast_1904_inst_req_1 : boolean;
  signal type_cast_1891_inst_ack_1 : boolean;
  signal type_cast_1891_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1900_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1918_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1918_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1869_inst_req_1 : boolean;
  signal type_cast_1904_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1860_inst_ack_1 : boolean;
  signal type_cast_1891_inst_ack_0 : boolean;
  signal type_cast_1963_inst_req_0 : boolean;
  signal type_cast_1963_inst_ack_0 : boolean;
  signal type_cast_1891_inst_req_0 : boolean;
  signal type_cast_1959_inst_req_1 : boolean;
  signal type_cast_1959_inst_ack_1 : boolean;
  signal type_cast_1959_inst_req_0 : boolean;
  signal type_cast_1959_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1887_inst_ack_1 : boolean;
  signal phi_stmt_1973_req_0 : boolean;
  signal RPIPE_Block1_start_1872_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1887_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1872_inst_req_1 : boolean;
  signal type_cast_1951_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1863_inst_ack_0 : boolean;
  signal type_cast_1963_inst_ack_1 : boolean;
  signal type_cast_1955_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1863_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1887_inst_ack_0 : boolean;
  signal type_cast_1963_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1887_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1872_inst_ack_0 : boolean;
  signal type_cast_1955_inst_req_0 : boolean;
  signal type_cast_2187_inst_ack_0 : boolean;
  signal type_cast_1955_inst_ack_0 : boolean;
  signal type_cast_1955_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1866_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1866_inst_req_1 : boolean;
  signal type_cast_1951_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1915_inst_req_1 : boolean;
  signal type_cast_1976_inst_ack_1 : boolean;
  signal type_cast_2034_inst_req_0 : boolean;
  signal type_cast_2034_inst_ack_0 : boolean;
  signal type_cast_2034_inst_req_1 : boolean;
  signal type_cast_2034_inst_ack_1 : boolean;
  signal type_cast_2038_inst_req_0 : boolean;
  signal type_cast_2038_inst_ack_0 : boolean;
  signal type_cast_2038_inst_req_1 : boolean;
  signal type_cast_2038_inst_ack_1 : boolean;
  signal type_cast_2042_inst_req_0 : boolean;
  signal type_cast_2042_inst_ack_0 : boolean;
  signal phi_stmt_2181_req_0 : boolean;
  signal type_cast_2042_inst_req_1 : boolean;
  signal type_cast_2042_inst_ack_1 : boolean;
  signal type_cast_2072_inst_req_0 : boolean;
  signal type_cast_2072_inst_ack_0 : boolean;
  signal type_cast_2072_inst_req_1 : boolean;
  signal type_cast_2072_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_0 : boolean;
  signal type_cast_2197_inst_ack_1 : boolean;
  signal array_obj_ref_2078_index_offset_req_0 : boolean;
  signal array_obj_ref_2078_index_offset_ack_0 : boolean;
  signal array_obj_ref_2078_index_offset_req_1 : boolean;
  signal array_obj_ref_2078_index_offset_ack_1 : boolean;
  signal type_cast_2197_inst_req_1 : boolean;
  signal addr_of_2079_final_reg_req_0 : boolean;
  signal addr_of_2079_final_reg_ack_0 : boolean;
  signal addr_of_2079_final_reg_req_1 : boolean;
  signal addr_of_2079_final_reg_ack_1 : boolean;
  signal type_cast_2197_inst_ack_0 : boolean;
  signal type_cast_2197_inst_req_0 : boolean;
  signal ptr_deref_2083_load_0_req_0 : boolean;
  signal ptr_deref_2083_load_0_ack_0 : boolean;
  signal ptr_deref_2083_load_0_req_1 : boolean;
  signal ptr_deref_2083_load_0_ack_1 : boolean;
  signal array_obj_ref_2101_index_offset_req_0 : boolean;
  signal array_obj_ref_2101_index_offset_ack_0 : boolean;
  signal array_obj_ref_2101_index_offset_req_1 : boolean;
  signal array_obj_ref_2101_index_offset_ack_1 : boolean;
  signal addr_of_2102_final_reg_req_0 : boolean;
  signal addr_of_2102_final_reg_ack_0 : boolean;
  signal addr_of_2102_final_reg_req_1 : boolean;
  signal addr_of_2102_final_reg_ack_1 : boolean;
  signal phi_stmt_2188_req_1 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_1 : boolean;
  signal ptr_deref_2105_store_0_req_0 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal ptr_deref_2105_store_0_ack_0 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal ptr_deref_2105_store_0_req_1 : boolean;
  signal ptr_deref_2105_store_0_ack_1 : boolean;
  signal type_cast_2110_inst_req_0 : boolean;
  signal type_cast_2110_inst_ack_0 : boolean;
  signal type_cast_2110_inst_req_1 : boolean;
  signal type_cast_2110_inst_ack_1 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal phi_stmt_2194_ack_0 : boolean;
  signal if_stmt_2123_branch_req_0 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal phi_stmt_2188_ack_0 : boolean;
  signal if_stmt_2123_branch_ack_1 : boolean;
  signal phi_stmt_2181_ack_0 : boolean;
  signal if_stmt_2123_branch_ack_0 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_2151_inst_req_0 : boolean;
  signal type_cast_2151_inst_ack_0 : boolean;
  signal type_cast_2151_inst_req_1 : boolean;
  signal type_cast_2151_inst_ack_1 : boolean;
  signal phi_stmt_2188_req_0 : boolean;
  signal type_cast_1976_inst_req_1 : boolean;
  signal type_cast_2167_inst_req_0 : boolean;
  signal type_cast_2167_inst_ack_0 : boolean;
  signal type_cast_2191_inst_ack_1 : boolean;
  signal type_cast_2167_inst_req_1 : boolean;
  signal type_cast_2167_inst_ack_1 : boolean;
  signal type_cast_2191_inst_req_1 : boolean;
  signal if_stmt_2174_branch_req_0 : boolean;
  signal phi_stmt_1994_ack_0 : boolean;
  signal if_stmt_2174_branch_ack_1 : boolean;
  signal if_stmt_2174_branch_ack_0 : boolean;
  signal phi_stmt_1987_ack_0 : boolean;
  signal phi_stmt_1980_ack_0 : boolean;
  signal type_cast_2191_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2210_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2210_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2210_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2210_inst_ack_1 : boolean;
  signal type_cast_2191_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_1999_inst_req_0 : boolean;
  signal type_cast_1999_inst_ack_0 : boolean;
  signal type_cast_1999_inst_req_1 : boolean;
  signal type_cast_1999_inst_ack_1 : boolean;
  signal phi_stmt_1994_req_1 : boolean;
  signal phi_stmt_1987_req_0 : boolean;
  signal phi_stmt_1980_req_0 : boolean;
  signal phi_stmt_1973_req_1 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_1997_inst_req_0 : boolean;
  signal type_cast_1997_inst_ack_0 : boolean;
  signal type_cast_1997_inst_req_1 : boolean;
  signal type_cast_1997_inst_ack_1 : boolean;
  signal phi_stmt_1994_req_0 : boolean;
  signal type_cast_1993_inst_req_0 : boolean;
  signal type_cast_1993_inst_ack_0 : boolean;
  signal type_cast_1993_inst_req_1 : boolean;
  signal type_cast_1993_inst_ack_1 : boolean;
  signal phi_stmt_1987_req_1 : boolean;
  signal type_cast_1986_inst_req_0 : boolean;
  signal type_cast_1986_inst_ack_0 : boolean;
  signal type_cast_1986_inst_req_1 : boolean;
  signal type_cast_1986_inst_ack_1 : boolean;
  signal phi_stmt_1980_req_1 : boolean;
  signal type_cast_1976_inst_req_0 : boolean;
  signal type_cast_1976_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4772_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4772_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4772_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4772_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4772: Block -- control-path 
    signal convTransposeB_CP_4772_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4772_elements(0) <= convTransposeB_CP_4772_start;
    convTransposeB_CP_4772_symbol <= convTransposeB_CP_4772_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1858/branch_block_stmt_1858__entry__
      -- CP-element group 0: 	 branch_block_stmt_1858/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919__entry__
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/$entry
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_sample_start_
      -- 
    rr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(0), ack => RPIPE_Block1_start_1860_inst_req_0); -- 
    cr_4993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(0), ack => type_cast_1904_inst_req_1); -- 
    cr_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(0), ack => type_cast_1891_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1858/assign_stmt_2206__exit__
      -- CP-element group 1: 	 branch_block_stmt_1858/assign_stmt_2206__entry__
      -- CP-element group 1: 	 branch_block_stmt_1858/merge_stmt_2180__exit__
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1858/assign_stmt_2206/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/assign_stmt_2206/$exit
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Sample/rr
      -- 
    cr_5595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1976_inst_req_1); -- 
    rr_5521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1997_inst_req_0); -- 
    cr_5526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1997_inst_req_1); -- 
    rr_5544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1993_inst_req_0); -- 
    cr_5549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1993_inst_req_1); -- 
    rr_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1986_inst_req_0); -- 
    cr_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1986_inst_req_1); -- 
    rr_5590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(1), ack => type_cast_1976_inst_req_0); -- 
    convTransposeB_CP_4772_elements(1) <= convTransposeB_CP_4772_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_sample_completed_
      -- 
    ra_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1860_inst_ack_0, ack => convTransposeB_CP_4772_elements(2)); -- 
    cr_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(2), ack => RPIPE_Block1_start_1860_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1860_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Sample/$entry
      -- 
    ca_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1860_inst_ack_1, ack => convTransposeB_CP_4772_elements(3)); -- 
    rr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(3), ack => RPIPE_Block1_start_1863_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_update_start_
      -- 
    ra_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1863_inst_ack_0, ack => convTransposeB_CP_4772_elements(4)); -- 
    cr_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(4), ack => RPIPE_Block1_start_1863_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1863_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_sample_start_
      -- 
    ca_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1863_inst_ack_1, ack => convTransposeB_CP_4772_elements(5)); -- 
    rr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(5), ack => RPIPE_Block1_start_1866_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Update/$entry
      -- 
    ra_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1866_inst_ack_0, ack => convTransposeB_CP_4772_elements(6)); -- 
    cr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(6), ack => RPIPE_Block1_start_1866_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1866_Update/$exit
      -- 
    ca_4854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1866_inst_ack_1, ack => convTransposeB_CP_4772_elements(7)); -- 
    rr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(7), ack => RPIPE_Block1_start_1869_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_sample_completed_
      -- 
    ra_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1869_inst_ack_0, ack => convTransposeB_CP_4772_elements(8)); -- 
    cr_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(8), ack => RPIPE_Block1_start_1869_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1869_Update/ca
      -- 
    ca_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1869_inst_ack_1, ack => convTransposeB_CP_4772_elements(9)); -- 
    rr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(9), ack => RPIPE_Block1_start_1872_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Sample/ra
      -- 
    ra_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1872_inst_ack_0, ack => convTransposeB_CP_4772_elements(10)); -- 
    cr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(10), ack => RPIPE_Block1_start_1872_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1872_Update/$exit
      -- 
    ca_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1872_inst_ack_1, ack => convTransposeB_CP_4772_elements(11)); -- 
    rr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(11), ack => RPIPE_Block1_start_1875_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_sample_completed_
      -- 
    ra_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1875_inst_ack_0, ack => convTransposeB_CP_4772_elements(12)); -- 
    cr_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(12), ack => RPIPE_Block1_start_1875_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1875_update_completed_
      -- 
    ca_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1875_inst_ack_1, ack => convTransposeB_CP_4772_elements(13)); -- 
    rr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(13), ack => RPIPE_Block1_start_1878_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Update/cr
      -- 
    ra_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1878_inst_ack_0, ack => convTransposeB_CP_4772_elements(14)); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(14), ack => RPIPE_Block1_start_1878_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1878_update_completed_
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1878_inst_ack_1, ack => convTransposeB_CP_4772_elements(15)); -- 
    rr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(15), ack => RPIPE_Block1_start_1881_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Sample/ra
      -- 
    ra_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1881_inst_ack_0, ack => convTransposeB_CP_4772_elements(16)); -- 
    cr_4923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(16), ack => RPIPE_Block1_start_1881_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1881_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_sample_start_
      -- 
    ca_4924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1881_inst_ack_1, ack => convTransposeB_CP_4772_elements(17)); -- 
    rr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(17), ack => RPIPE_Block1_start_1884_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_sample_completed_
      -- 
    ra_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1884_inst_ack_0, ack => convTransposeB_CP_4772_elements(18)); -- 
    cr_4937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(18), ack => RPIPE_Block1_start_1884_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1884_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Sample/rr
      -- 
    ca_4938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1884_inst_ack_1, ack => convTransposeB_CP_4772_elements(19)); -- 
    rr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(19), ack => RPIPE_Block1_start_1887_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Sample/ra
      -- 
    ra_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1887_inst_ack_0, ack => convTransposeB_CP_4772_elements(20)); -- 
    cr_4951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(20), ack => RPIPE_Block1_start_1887_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1887_Update/$exit
      -- 
    ca_4952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1887_inst_ack_1, ack => convTransposeB_CP_4772_elements(21)); -- 
    rr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(21), ack => type_cast_1891_inst_req_0); -- 
    rr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(21), ack => RPIPE_Block1_start_1900_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_sample_completed_
      -- 
    ra_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1891_inst_ack_0, ack => convTransposeB_CP_4772_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1891_update_completed_
      -- 
    ca_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1891_inst_ack_1, ack => convTransposeB_CP_4772_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Update/cr
      -- 
    ra_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1900_inst_ack_0, ack => convTransposeB_CP_4772_elements(24)); -- 
    cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(24), ack => RPIPE_Block1_start_1900_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1900_Update/ca
      -- 
    ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1900_inst_ack_1, ack => convTransposeB_CP_4772_elements(25)); -- 
    rr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(25), ack => type_cast_1904_inst_req_0); -- 
    rr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(25), ack => RPIPE_Block1_start_1912_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Sample/$exit
      -- 
    ra_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1904_inst_ack_0, ack => convTransposeB_CP_4772_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/type_cast_1904_Update/ca
      -- 
    ca_4994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1904_inst_ack_1, ack => convTransposeB_CP_4772_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Sample/$exit
      -- 
    ra_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1912_inst_ack_0, ack => convTransposeB_CP_4772_elements(28)); -- 
    cr_5007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(28), ack => RPIPE_Block1_start_1912_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1912_update_completed_
      -- 
    ca_5008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1912_inst_ack_1, ack => convTransposeB_CP_4772_elements(29)); -- 
    rr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(29), ack => RPIPE_Block1_start_1915_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Update/cr
      -- 
    ra_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1915_inst_ack_0, ack => convTransposeB_CP_4772_elements(30)); -- 
    cr_5021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(30), ack => RPIPE_Block1_start_1915_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1915_Update/$exit
      -- 
    ca_5022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1915_inst_ack_1, ack => convTransposeB_CP_4772_elements(31)); -- 
    rr_5030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(31), ack => RPIPE_Block1_start_1918_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Sample/ra
      -- 
    ra_5031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1918_inst_ack_0, ack => convTransposeB_CP_4772_elements(32)); -- 
    cr_5035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(32), ack => RPIPE_Block1_start_1918_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/RPIPE_Block1_start_1918_update_completed_
      -- 
    ca_5036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1918_inst_ack_1, ack => convTransposeB_CP_4772_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970__entry__
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919__exit__
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1861_to_assign_stmt_1919/$exit
      -- CP-element group 34: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Sample/$entry
      -- 
    rr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1951_inst_req_0); -- 
    rr_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1963_inst_req_0); -- 
    cr_5080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1959_inst_req_1); -- 
    rr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1959_inst_req_0); -- 
    cr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1951_inst_req_1); -- 
    cr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1955_inst_req_1); -- 
    cr_5094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1963_inst_req_1); -- 
    rr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(34), ack => type_cast_1955_inst_req_0); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(23) & convTransposeB_CP_4772_elements(27) & convTransposeB_CP_4772_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Sample/$exit
      -- 
    ra_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_0, ack => convTransposeB_CP_4772_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1951_update_completed_
      -- 
    ca_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_1, ack => convTransposeB_CP_4772_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_sample_completed_
      -- 
    ra_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_0, ack => convTransposeB_CP_4772_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1955_update_completed_
      -- 
    ca_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_1, ack => convTransposeB_CP_4772_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_sample_completed_
      -- 
    ra_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1959_inst_ack_0, ack => convTransposeB_CP_4772_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1959_update_completed_
      -- 
    ca_5081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1959_inst_ack_1, ack => convTransposeB_CP_4772_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_sample_completed_
      -- 
    ra_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1963_inst_ack_0, ack => convTransposeB_CP_4772_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/type_cast_1963_Update/$exit
      -- 
    ca_5095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1963_inst_ack_1, ack => convTransposeB_CP_4772_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970__exit__
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1858/assign_stmt_1926_to_assign_stmt_1970/$exit
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1987/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1980/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1973/$entry
      -- CP-element group 43: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$entry
      -- 
    rr_5471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(43), ack => type_cast_1999_inst_req_0); -- 
    cr_5476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(43), ack => type_cast_1999_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(36) & convTransposeB_CP_4772_elements(38) & convTransposeB_CP_4772_elements(40) & convTransposeB_CP_4772_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Sample/ra
      -- 
    ra_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2034_inst_ack_0, ack => convTransposeB_CP_4772_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Update/ca
      -- 
    ca_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2034_inst_ack_1, ack => convTransposeB_CP_4772_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Sample/ra
      -- 
    ra_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_0, ack => convTransposeB_CP_4772_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Update/ca
      -- 
    ca_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_1, ack => convTransposeB_CP_4772_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Sample/ra
      -- 
    ra_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2042_inst_ack_0, ack => convTransposeB_CP_4772_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Update/ca
      -- 
    ca_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2042_inst_ack_1, ack => convTransposeB_CP_4772_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Sample/ra
      -- 
    ra_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2072_inst_ack_0, ack => convTransposeB_CP_4772_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Sample/req
      -- 
    ca_5154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2072_inst_ack_1, ack => convTransposeB_CP_4772_elements(51)); -- 
    req_5179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(51), ack => array_obj_ref_2078_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Sample/ack
      -- 
    ack_5180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2078_index_offset_ack_0, ack => convTransposeB_CP_4772_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_request/req
      -- 
    ack_5185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2078_index_offset_ack_1, ack => convTransposeB_CP_4772_elements(53)); -- 
    req_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(53), ack => addr_of_2079_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_request/ack
      -- 
    ack_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2079_final_reg_ack_0, ack => convTransposeB_CP_4772_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/word_access_start/word_0/rr
      -- 
    ack_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2079_final_reg_ack_1, ack => convTransposeB_CP_4772_elements(55)); -- 
    rr_5233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(55), ack => ptr_deref_2083_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Sample/word_access_start/word_0/ra
      -- 
    ra_5234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2083_load_0_ack_0, ack => convTransposeB_CP_4772_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/ptr_deref_2083_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/ptr_deref_2083_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/ptr_deref_2083_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/ptr_deref_2083_Merge/merge_ack
      -- 
    ca_5245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2083_load_0_ack_1, ack => convTransposeB_CP_4772_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Sample/req
      -- 
    req_5275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(58), ack => array_obj_ref_2101_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(45) & convTransposeB_CP_4772_elements(47) & convTransposeB_CP_4772_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Sample/ack
      -- 
    ack_5276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2101_index_offset_ack_0, ack => convTransposeB_CP_4772_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_request/req
      -- 
    ack_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2101_index_offset_ack_1, ack => convTransposeB_CP_4772_elements(60)); -- 
    req_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(60), ack => addr_of_2102_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_request/ack
      -- 
    ack_5291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2102_final_reg_ack_0, ack => convTransposeB_CP_4772_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_word_addrgen/root_register_ack
      -- 
    ack_5296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2102_final_reg_ack_1, ack => convTransposeB_CP_4772_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/ptr_deref_2105_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/ptr_deref_2105_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/ptr_deref_2105_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/ptr_deref_2105_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/word_access_start/word_0/rr
      -- 
    rr_5334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(63), ack => ptr_deref_2105_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(57) & convTransposeB_CP_4772_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Sample/word_access_start/word_0/ra
      -- 
    ra_5335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2105_store_0_ack_0, ack => convTransposeB_CP_4772_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/word_access_complete/word_0/ca
      -- 
    ca_5346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2105_store_0_ack_1, ack => convTransposeB_CP_4772_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Sample/ra
      -- 
    ra_5355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2110_inst_ack_0, ack => convTransposeB_CP_4772_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Update/ca
      -- 
    ca_5360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2110_inst_ack_1, ack => convTransposeB_CP_4772_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122__exit__
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123__entry__
      -- CP-element group 68: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/$exit
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1858/R_cmp_2124_place
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1858/if_stmt_2123_else_link/$entry
      -- 
    branch_req_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(68), ack => if_stmt_2123_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(52) & convTransposeB_CP_4772_elements(59) & convTransposeB_CP_4772_elements(65) & convTransposeB_CP_4772_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/assign_stmt_2135__entry__
      -- CP-element group 69: 	 branch_block_stmt_1858/assign_stmt_2135__exit__
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1858/merge_stmt_2129__exit__
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/merge_stmt_2129_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1858/merge_stmt_2129_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1858/merge_stmt_2129_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1858/if_stmt_2123_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1858/merge_stmt_2129_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/if_stmt_2123_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1858/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1858/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1858/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/assign_stmt_2135/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/assign_stmt_2135/$exit
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/rr
      -- 
    if_choice_transition_5373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2123_branch_ack_1, ack => convTransposeB_CP_4772_elements(69)); -- 
    cr_5733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2187_inst_req_1); -- 
    rr_5728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2187_inst_req_0); -- 
    cr_5710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2197_inst_req_1); -- 
    rr_5705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2197_inst_req_0); -- 
    cr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2191_inst_req_1); -- 
    rr_5751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(69), ack => type_cast_2191_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173__entry__
      -- CP-element group 70: 	 branch_block_stmt_1858/merge_stmt_2137__exit__
      -- CP-element group 70: 	 branch_block_stmt_1858/merge_stmt_2137_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1858/merge_stmt_2137_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1858/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1858/merge_stmt_2137_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1858/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1858/if_stmt_2123_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1858/if_stmt_2123_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1858/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/$entry
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1858/merge_stmt_2137_PhiAck/dummy
      -- 
    else_choice_transition_5377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2123_branch_ack_0, ack => convTransposeB_CP_4772_elements(70)); -- 
    rr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(70), ack => type_cast_2151_inst_req_0); -- 
    cr_5398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(70), ack => type_cast_2151_inst_req_1); -- 
    cr_5412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(70), ack => type_cast_2167_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Sample/ra
      -- 
    ra_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2151_inst_ack_0, ack => convTransposeB_CP_4772_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2151_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Sample/rr
      -- 
    ca_5399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2151_inst_ack_1, ack => convTransposeB_CP_4772_elements(72)); -- 
    rr_5407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(72), ack => type_cast_2167_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Sample/ra
      -- 
    ra_5408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2167_inst_ack_0, ack => convTransposeB_CP_4772_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174__entry__
      -- CP-element group 74: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173__exit__
      -- CP-element group 74: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/$exit
      -- CP-element group 74: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1858/assign_stmt_2143_to_assign_stmt_2173/type_cast_2167_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1858/R_cmp117_2175_place
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1858/if_stmt_2174_else_link/$entry
      -- 
    ca_5413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2167_inst_ack_1, ack => convTransposeB_CP_4772_elements(74)); -- 
    branch_req_5421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(74), ack => if_stmt_2174_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1858/merge_stmt_2208__exit__
      -- CP-element group 75: 	 branch_block_stmt_1858/assign_stmt_2213__entry__
      -- CP-element group 75: 	 branch_block_stmt_1858/merge_stmt_2208_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1858/merge_stmt_2208_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1858/merge_stmt_2208_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1858/merge_stmt_2208_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1858/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1858/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1858/if_stmt_2174_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1858/if_stmt_2174_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1858/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1858/assign_stmt_2213/$entry
      -- CP-element group 75: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Sample/req
      -- 
    if_choice_transition_5426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2174_branch_ack_1, ack => convTransposeB_CP_4772_elements(75)); -- 
    req_5446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(75), ack => WPIPE_Block1_done_2210_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2181/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/if_stmt_2174_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1858/if_stmt_2174_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/$entry
      -- CP-element group 76: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$entry
      -- 
    else_choice_transition_5430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2174_branch_ack_0, ack => convTransposeB_CP_4772_elements(76)); -- 
    cr_5684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2193_inst_req_1); -- 
    rr_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2193_inst_req_0); -- 
    cr_5653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2199_inst_req_1); -- 
    rr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(76), ack => type_cast_2199_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Update/req
      -- 
    ack_5447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2210_inst_ack_0, ack => convTransposeB_CP_4772_elements(77)); -- 
    req_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(77), ack => WPIPE_Block1_done_2210_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1858/$exit
      -- CP-element group 78: 	 branch_block_stmt_1858/return__
      -- CP-element group 78: 	 branch_block_stmt_1858/branch_block_stmt_1858__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1858/merge_stmt_2215__exit__
      -- CP-element group 78: 	 branch_block_stmt_1858/assign_stmt_2213__exit__
      -- CP-element group 78: 	 branch_block_stmt_1858/merge_stmt_2215_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1858/merge_stmt_2215_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1858/merge_stmt_2215_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1858/merge_stmt_2215_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1858/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1858/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1858/assign_stmt_2213/$exit
      -- CP-element group 78: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1858/assign_stmt_2213/WPIPE_Block1_done_2210_Update/ack
      -- 
    ack_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2210_inst_ack_1, ack => convTransposeB_CP_4772_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Sample/ra
      -- 
    ra_5472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_0, ack => convTransposeB_CP_4772_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/Update/ca
      -- 
    ca_5477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_1, ack => convTransposeB_CP_4772_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/$exit
      -- CP-element group 81: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/$exit
      -- CP-element group 81: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1999/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_req
      -- 
    phi_stmt_1994_req_5478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1994_req_5478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(81), ack => phi_stmt_1994_req_1); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(79) & convTransposeB_CP_4772_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1987/$exit
      -- CP-element group 82: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1991_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_req
      -- 
    phi_stmt_1987_req_5486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1987_req_5486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(82), ack => phi_stmt_1987_req_0); -- 
    -- Element group convTransposeB_CP_4772_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(43), ack => convTransposeB_CP_4772_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1980/$exit
      -- CP-element group 83: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1984_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_req
      -- 
    phi_stmt_1980_req_5494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1980_req_5494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(83), ack => phi_stmt_1980_req_0); -- 
    -- Element group convTransposeB_CP_4772_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(43), ack => convTransposeB_CP_4772_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1973/$exit
      -- CP-element group 84: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_req
      -- 
    phi_stmt_1973_req_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1973_req_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(84), ack => phi_stmt_1973_req_1); -- 
    -- Element group convTransposeB_CP_4772_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(43), ack => convTransposeB_CP_4772_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1858/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(81) & convTransposeB_CP_4772_elements(82) & convTransposeB_CP_4772_elements(83) & convTransposeB_CP_4772_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Sample/ra
      -- 
    ra_5522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1997_inst_ack_0, ack => convTransposeB_CP_4772_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/Update/ca
      -- 
    ca_5527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1997_inst_ack_1, ack => convTransposeB_CP_4772_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/$exit
      -- CP-element group 88: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/$exit
      -- CP-element group 88: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_sources/type_cast_1997/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1994/phi_stmt_1994_req
      -- 
    phi_stmt_1994_req_5528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1994_req_5528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(88), ack => phi_stmt_1994_req_0); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(86) & convTransposeB_CP_4772_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Sample/ra
      -- 
    ra_5545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_0, ack => convTransposeB_CP_4772_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/Update/ca
      -- 
    ca_5550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_1, ack => convTransposeB_CP_4772_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/$exit
      -- CP-element group 91: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/$exit
      -- CP-element group 91: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_sources/type_cast_1993/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1987/phi_stmt_1987_req
      -- 
    phi_stmt_1987_req_5551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1987_req_5551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(91), ack => phi_stmt_1987_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(89) & convTransposeB_CP_4772_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Sample/ra
      -- 
    ra_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1986_inst_ack_0, ack => convTransposeB_CP_4772_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/Update/ca
      -- 
    ca_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1986_inst_ack_1, ack => convTransposeB_CP_4772_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/$exit
      -- CP-element group 94: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/$exit
      -- CP-element group 94: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_sources/type_cast_1986/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1980/phi_stmt_1980_req
      -- 
    phi_stmt_1980_req_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1980_req_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(94), ack => phi_stmt_1980_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(92) & convTransposeB_CP_4772_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Sample/ra
      -- 
    ra_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_0, ack => convTransposeB_CP_4772_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/Update/$exit
      -- 
    ca_5596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_1, ack => convTransposeB_CP_4772_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_req
      -- CP-element group 97: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/$exit
      -- CP-element group 97: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/$exit
      -- CP-element group 97: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1976/SplitProtocol/$exit
      -- 
    phi_stmt_1973_req_5597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1973_req_5597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(97), ack => phi_stmt_1973_req_0); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(95) & convTransposeB_CP_4772_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1858/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(88) & convTransposeB_CP_4772_elements(91) & convTransposeB_CP_4772_elements(94) & convTransposeB_CP_4772_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1858/merge_stmt_1972_PhiAck/$entry
      -- CP-element group 99: 	 branch_block_stmt_1858/merge_stmt_1972_PhiReqMerge
      -- 
    convTransposeB_CP_4772_elements(99) <= OrReduce(convTransposeB_CP_4772_elements(85) & convTransposeB_CP_4772_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1858/merge_stmt_1972_PhiAck/phi_stmt_1973_ack
      -- 
    phi_stmt_1973_ack_5602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1973_ack_0, ack => convTransposeB_CP_4772_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1858/merge_stmt_1972_PhiAck/phi_stmt_1980_ack
      -- 
    phi_stmt_1980_ack_5603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1980_ack_0, ack => convTransposeB_CP_4772_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1858/merge_stmt_1972_PhiAck/phi_stmt_1987_ack
      -- 
    phi_stmt_1987_ack_5604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1987_ack_0, ack => convTransposeB_CP_4772_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1858/merge_stmt_1972_PhiAck/phi_stmt_1994_ack
      -- 
    phi_stmt_1994_ack_5605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1994_ack_0, ack => convTransposeB_CP_4772_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122__entry__
      -- CP-element group 104: 	 branch_block_stmt_1858/merge_stmt_1972_PhiAck/$exit
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/merge_stmt_1972__exit__
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2034_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2038_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2042_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2072_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2078_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2079_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2083_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/array_obj_ref_2101_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/addr_of_2102_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/ptr_deref_2105_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1858/assign_stmt_2006_to_assign_stmt_2122/type_cast_2110_Update/cr
      -- 
    rr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2034_inst_req_0); -- 
    cr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2034_inst_req_1); -- 
    rr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2038_inst_req_0); -- 
    cr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2038_inst_req_1); -- 
    rr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2042_inst_req_0); -- 
    cr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2042_inst_req_1); -- 
    rr_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2072_inst_req_0); -- 
    cr_5153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2072_inst_req_1); -- 
    req_5184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => array_obj_ref_2078_index_offset_req_1); -- 
    req_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => addr_of_2079_final_reg_req_1); -- 
    cr_5244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => ptr_deref_2083_load_0_req_1); -- 
    req_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => array_obj_ref_2101_index_offset_req_1); -- 
    req_5295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => addr_of_2102_final_reg_req_1); -- 
    cr_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => ptr_deref_2105_store_0_req_1); -- 
    rr_5354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2110_inst_req_0); -- 
    cr_5359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(104), ack => type_cast_2110_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(100) & convTransposeB_CP_4772_elements(101) & convTransposeB_CP_4772_elements(102) & convTransposeB_CP_4772_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$exit
      -- 
    ra_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => convTransposeB_CP_4772_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$exit
      -- 
    ca_5654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => convTransposeB_CP_4772_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$exit
      -- CP-element group 107: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/$exit
      -- CP-element group 107: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    phi_stmt_2194_req_5655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2194_req_5655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(107), ack => phi_stmt_2194_req_1); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(105) & convTransposeB_CP_4772_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_req
      -- CP-element group 108: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2185_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2181/$exit
      -- 
    phi_stmt_2181_req_5663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2181_req_5663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(108), ack => phi_stmt_2181_req_0); -- 
    -- Element group convTransposeB_CP_4772_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => convTransposeB_CP_4772_elements(76), ack => convTransposeB_CP_4772_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- 
    ra_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => convTransposeB_CP_4772_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/ca
      -- CP-element group 110: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- 
    ca_5685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => convTransposeB_CP_4772_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/$exit
      -- CP-element group 111: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_req
      -- CP-element group 111: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2193/$exit
      -- CP-element group 111: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$exit
      -- 
    phi_stmt_2188_req_5686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2188_req_5686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(111), ack => phi_stmt_2188_req_1); -- 
    convTransposeB_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(109) & convTransposeB_CP_4772_elements(110);
      gj_convTransposeB_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1858/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(107) & convTransposeB_CP_4772_elements(108) & convTransposeB_CP_4772_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$exit
      -- 
    ra_5706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_0, ack => convTransposeB_CP_4772_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$exit
      -- 
    ca_5711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_1, ack => convTransposeB_CP_4772_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- CP-element group 115: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$exit
      -- CP-element group 115: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2194/$exit
      -- 
    phi_stmt_2194_req_5712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2194_req_5712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(115), ack => phi_stmt_2194_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(113) & convTransposeB_CP_4772_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Sample/ra
      -- 
    ra_5729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_0, ack => convTransposeB_CP_4772_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/Update/$exit
      -- 
    ca_5734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_1, ack => convTransposeB_CP_4772_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_req
      -- CP-element group 118: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2187/$exit
      -- CP-element group 118: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2181/$exit
      -- 
    phi_stmt_2181_req_5735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2181_req_5735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(118), ack => phi_stmt_2181_req_1); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(116) & convTransposeB_CP_4772_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Sample/$exit
      -- 
    ra_5752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2191_inst_ack_0, ack => convTransposeB_CP_4772_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/Update/$exit
      -- 
    ca_5757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2191_inst_ack_1, ack => convTransposeB_CP_4772_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/$exit
      -- CP-element group 121: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_sources/type_cast_2191/$exit
      -- CP-element group 121: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2188/phi_stmt_2188_req
      -- 
    phi_stmt_2188_req_5758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2188_req_5758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4772_elements(121), ack => phi_stmt_2188_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(119) & convTransposeB_CP_4772_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1858/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(115) & convTransposeB_CP_4772_elements(118) & convTransposeB_CP_4772_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1858/merge_stmt_2180_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1858/merge_stmt_2180_PhiAck/$entry
      -- 
    convTransposeB_CP_4772_elements(123) <= OrReduce(convTransposeB_CP_4772_elements(112) & convTransposeB_CP_4772_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1858/merge_stmt_2180_PhiAck/phi_stmt_2181_ack
      -- 
    phi_stmt_2181_ack_5763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2181_ack_0, ack => convTransposeB_CP_4772_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1858/merge_stmt_2180_PhiAck/phi_stmt_2188_ack
      -- 
    phi_stmt_2188_ack_5764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2188_ack_0, ack => convTransposeB_CP_4772_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1858/merge_stmt_2180_PhiAck/phi_stmt_2194_ack
      -- 
    phi_stmt_2194_ack_5765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2194_ack_0, ack => convTransposeB_CP_4772_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1858/merge_stmt_2180_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4772_elements(124) & convTransposeB_CP_4772_elements(125) & convTransposeB_CP_4772_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4772_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2100_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2100_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2077_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2077_scaled : std_logic_vector(13 downto 0);
    signal add45_1932 : std_logic_vector(15 downto 0);
    signal add58_1943 : std_logic_vector(15 downto 0);
    signal add77_2053 : std_logic_vector(63 downto 0);
    signal add79_2063 : std_logic_vector(63 downto 0);
    signal add91_2117 : std_logic_vector(31 downto 0);
    signal add98_2135 : std_logic_vector(15 downto 0);
    signal add_1910 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2011 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2078_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2078_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2078_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2078_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2078_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2078_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2101_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2101_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2101_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2101_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2101_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2101_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2080 : std_logic_vector(31 downto 0);
    signal arrayidx87_2103 : std_logic_vector(31 downto 0);
    signal call11_1879 : std_logic_vector(15 downto 0);
    signal call13_1882 : std_logic_vector(15 downto 0);
    signal call14_1885 : std_logic_vector(15 downto 0);
    signal call15_1888 : std_logic_vector(15 downto 0);
    signal call16_1901 : std_logic_vector(15 downto 0);
    signal call18_1913 : std_logic_vector(15 downto 0);
    signal call1_1864 : std_logic_vector(15 downto 0);
    signal call20_1916 : std_logic_vector(15 downto 0);
    signal call22_1919 : std_logic_vector(15 downto 0);
    signal call3_1867 : std_logic_vector(15 downto 0);
    signal call5_1870 : std_logic_vector(15 downto 0);
    signal call7_1873 : std_logic_vector(15 downto 0);
    signal call9_1876 : std_logic_vector(15 downto 0);
    signal call_1861 : std_logic_vector(15 downto 0);
    signal cmp106_2148 : std_logic_vector(0 downto 0);
    signal cmp117_2173 : std_logic_vector(0 downto 0);
    signal cmp_2122 : std_logic_vector(0 downto 0);
    signal conv112_2168 : std_logic_vector(31 downto 0);
    signal conv115_1964 : std_logic_vector(31 downto 0);
    signal conv17_1905 : std_logic_vector(31 downto 0);
    signal conv65_2035 : std_logic_vector(63 downto 0);
    signal conv68_1952 : std_logic_vector(63 downto 0);
    signal conv70_2039 : std_logic_vector(63 downto 0);
    signal conv73_1956 : std_logic_vector(63 downto 0);
    signal conv75_2043 : std_logic_vector(63 downto 0);
    signal conv90_2111 : std_logic_vector(31 downto 0);
    signal conv94_1960 : std_logic_vector(31 downto 0);
    signal conv_1892 : std_logic_vector(31 downto 0);
    signal idxprom86_2096 : std_logic_vector(63 downto 0);
    signal idxprom_2073 : std_logic_vector(63 downto 0);
    signal inc110_2152 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2157 : std_logic_vector(15 downto 0);
    signal inc_2143 : std_logic_vector(15 downto 0);
    signal indvar_1973 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2206 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2194 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1994 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2188 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1987 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2164 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2181 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1980 : std_logic_vector(15 downto 0);
    signal mul54_2026 : std_logic_vector(15 downto 0);
    signal mul76_2048 : std_logic_vector(63 downto 0);
    signal mul78_2058 : std_logic_vector(63 downto 0);
    signal mul_2016 : std_logic_vector(15 downto 0);
    signal ptr_deref_2083_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2083_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2083_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2083_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2083_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2105_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2105_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2105_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2105_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2105_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2105_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1898 : std_logic_vector(31 downto 0);
    signal shr116132_1970 : std_logic_vector(31 downto 0);
    signal shr131_1926 : std_logic_vector(15 downto 0);
    signal shr81_2069 : std_logic_vector(31 downto 0);
    signal shr85_2090 : std_logic_vector(63 downto 0);
    signal sub48_2021 : std_logic_vector(15 downto 0);
    signal sub61_1948 : std_logic_vector(15 downto 0);
    signal sub62_2031 : std_logic_vector(15 downto 0);
    signal sub_1937 : std_logic_vector(15 downto 0);
    signal tmp1_2006 : std_logic_vector(31 downto 0);
    signal tmp83_2084 : std_logic_vector(63 downto 0);
    signal type_cast_1896_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1924_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1930_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1941_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1968_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1976_wire : std_logic_vector(31 downto 0);
    signal type_cast_1979_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1984_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1986_wire : std_logic_vector(15 downto 0);
    signal type_cast_1991_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1993_wire : std_logic_vector(15 downto 0);
    signal type_cast_1997_wire : std_logic_vector(15 downto 0);
    signal type_cast_1999_wire : std_logic_vector(15 downto 0);
    signal type_cast_2004_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2067_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2088_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2094_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2115_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2133_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2141_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2161_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2185_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2187_wire : std_logic_vector(15 downto 0);
    signal type_cast_2191_wire : std_logic_vector(15 downto 0);
    signal type_cast_2193_wire : std_logic_vector(15 downto 0);
    signal type_cast_2197_wire : std_logic_vector(15 downto 0);
    signal type_cast_2199_wire : std_logic_vector(15 downto 0);
    signal type_cast_2204_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2212_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2078_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2078_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2078_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2078_resized_base_address <= "00000000000000";
    array_obj_ref_2101_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2101_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2101_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2101_resized_base_address <= "00000000000000";
    ptr_deref_2083_word_offset_0 <= "00000000000000";
    ptr_deref_2105_word_offset_0 <= "00000000000000";
    type_cast_1896_wire_constant <= "00000000000000000000000000010000";
    type_cast_1924_wire_constant <= "0000000000000010";
    type_cast_1930_wire_constant <= "1111111111111111";
    type_cast_1941_wire_constant <= "1111111111111111";
    type_cast_1968_wire_constant <= "00000000000000000000000000000001";
    type_cast_1979_wire_constant <= "00000000000000000000000000000000";
    type_cast_1984_wire_constant <= "0000000000000000";
    type_cast_1991_wire_constant <= "0000000000000000";
    type_cast_2004_wire_constant <= "00000000000000000000000000000100";
    type_cast_2067_wire_constant <= "00000000000000000000000000000010";
    type_cast_2088_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2094_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2115_wire_constant <= "00000000000000000000000000000100";
    type_cast_2133_wire_constant <= "0000000000000100";
    type_cast_2141_wire_constant <= "0000000000000001";
    type_cast_2161_wire_constant <= "0000000000000000";
    type_cast_2185_wire_constant <= "0000000000000000";
    type_cast_2204_wire_constant <= "00000000000000000000000000000001";
    type_cast_2212_wire_constant <= "0000000000000001";
    phi_stmt_1973: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1976_wire & type_cast_1979_wire_constant;
      req <= phi_stmt_1973_req_0 & phi_stmt_1973_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1973",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1973_ack_0,
          idata => idata,
          odata => indvar_1973,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1973
    phi_stmt_1980: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1984_wire_constant & type_cast_1986_wire;
      req <= phi_stmt_1980_req_0 & phi_stmt_1980_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1980",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1980_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1980,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1980
    phi_stmt_1987: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1991_wire_constant & type_cast_1993_wire;
      req <= phi_stmt_1987_req_0 & phi_stmt_1987_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1987",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1987_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1987,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1987
    phi_stmt_1994: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1997_wire & type_cast_1999_wire;
      req <= phi_stmt_1994_req_0 & phi_stmt_1994_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1994",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1994_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1994,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1994
    phi_stmt_2181: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2185_wire_constant & type_cast_2187_wire;
      req <= phi_stmt_2181_req_0 & phi_stmt_2181_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2181",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2181_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2181,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2181
    phi_stmt_2188: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2191_wire & type_cast_2193_wire;
      req <= phi_stmt_2188_req_0 & phi_stmt_2188_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2188",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2188_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2188,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2188
    phi_stmt_2194: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2197_wire & type_cast_2199_wire;
      req <= phi_stmt_2194_req_0 & phi_stmt_2194_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2194",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2194_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2194,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2194
    -- flow-through select operator MUX_2163_inst
    input_dim1x_x2_2164 <= type_cast_2161_wire_constant when (cmp106_2148(0) /=  '0') else inc_2143;
    addr_of_2079_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2079_final_reg_req_0;
      addr_of_2079_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2079_final_reg_req_1;
      addr_of_2079_final_reg_ack_1<= rack(0);
      addr_of_2079_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2079_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2078_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2080,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2102_final_reg_req_0;
      addr_of_2102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2102_final_reg_req_1;
      addr_of_2102_final_reg_ack_1<= rack(0);
      addr_of_2102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1891_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1891_inst_req_0;
      type_cast_1891_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1891_inst_req_1;
      type_cast_1891_inst_ack_1<= rack(0);
      type_cast_1891_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1891_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1888,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1892,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1904_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1904_inst_req_0;
      type_cast_1904_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1904_inst_req_1;
      type_cast_1904_inst_ack_1<= rack(0);
      type_cast_1904_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1904_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1905,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1951_inst_req_0;
      type_cast_1951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1951_inst_req_1;
      type_cast_1951_inst_ack_1<= rack(0);
      type_cast_1951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1919,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1955_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1955_inst_req_0;
      type_cast_1955_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1955_inst_req_1;
      type_cast_1955_inst_ack_1<= rack(0);
      type_cast_1955_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1955_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1959_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1959_inst_req_0;
      type_cast_1959_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1959_inst_req_1;
      type_cast_1959_inst_ack_1<= rack(0);
      type_cast_1959_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1959_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1960,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1963_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1963_inst_req_0;
      type_cast_1963_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1963_inst_req_1;
      type_cast_1963_inst_ack_1<= rack(0);
      type_cast_1963_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1963_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1964,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1976_inst_req_0;
      type_cast_1976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1976_inst_req_1;
      type_cast_1976_inst_ack_1<= rack(0);
      type_cast_1976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2206,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1976_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1986_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1986_inst_req_0;
      type_cast_1986_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1986_inst_req_1;
      type_cast_1986_inst_ack_1<= rack(0);
      type_cast_1986_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1986_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1986_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1993_inst_req_0;
      type_cast_1993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1993_inst_req_1;
      type_cast_1993_inst_ack_1<= rack(0);
      type_cast_1993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1993_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1997_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1997_inst_req_0;
      type_cast_1997_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1997_inst_req_1;
      type_cast_1997_inst_ack_1<= rack(0);
      type_cast_1997_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1997_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1997_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1999_inst_req_0;
      type_cast_1999_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1999_inst_req_1;
      type_cast_1999_inst_ack_1<= rack(0);
      type_cast_1999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1999_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1999_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2034_inst_req_0;
      type_cast_2034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2034_inst_req_1;
      type_cast_2034_inst_ack_1<= rack(0);
      type_cast_2034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1980,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2038_inst_req_0;
      type_cast_2038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2038_inst_req_1;
      type_cast_2038_inst_ack_1<= rack(0);
      type_cast_2038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2031,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2042_inst_req_0;
      type_cast_2042_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2042_inst_req_1;
      type_cast_2042_inst_ack_1<= rack(0);
      type_cast_2042_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2042_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2021,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2043,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2072_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2072_inst_req_0;
      type_cast_2072_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2072_inst_req_1;
      type_cast_2072_inst_ack_1<= rack(0);
      type_cast_2072_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2072_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2069,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2073,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2110_inst_req_0;
      type_cast_2110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2110_inst_req_1;
      type_cast_2110_inst_ack_1<= rack(0);
      type_cast_2110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1980,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2151_inst_req_0;
      type_cast_2151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2151_inst_req_1;
      type_cast_2151_inst_ack_1<= rack(0);
      type_cast_2151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2167_inst_req_0;
      type_cast_2167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2167_inst_req_1;
      type_cast_2167_inst_ack_1<= rack(0);
      type_cast_2167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2187_inst_req_0;
      type_cast_2187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2187_inst_req_1;
      type_cast_2187_inst_ack_1<= rack(0);
      type_cast_2187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2187_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2191_inst_req_0;
      type_cast_2191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2191_inst_req_1;
      type_cast_2191_inst_ack_1<= rack(0);
      type_cast_2191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1987,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2191_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2164,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2197_inst_req_0;
      type_cast_2197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2197_inst_req_1;
      type_cast_2197_inst_ack_1<= rack(0);
      type_cast_2197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1994,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2197_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2199_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2078_index_1_rename
    process(R_idxprom_2077_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2077_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2077_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2078_index_1_resize
    process(idxprom_2073) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2073;
      ov := iv(13 downto 0);
      R_idxprom_2077_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2078_root_address_inst
    process(array_obj_ref_2078_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2078_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2078_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2101_index_1_rename
    process(R_idxprom86_2100_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2100_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2100_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2101_index_1_resize
    process(idxprom86_2096) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2096;
      ov := iv(13 downto 0);
      R_idxprom86_2100_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2101_root_address_inst
    process(array_obj_ref_2101_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2101_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2101_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_addr_0
    process(ptr_deref_2083_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2083_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2083_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_base_resize
    process(arrayidx82_2080) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2080;
      ov := iv(13 downto 0);
      ptr_deref_2083_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_gather_scatter
    process(ptr_deref_2083_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2083_data_0;
      ov(63 downto 0) := iv;
      tmp83_2084 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_root_address_inst
    process(ptr_deref_2083_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2083_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2083_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2105_addr_0
    process(ptr_deref_2105_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2105_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2105_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2105_base_resize
    process(arrayidx87_2103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2103;
      ov := iv(13 downto 0);
      ptr_deref_2105_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2105_gather_scatter
    process(tmp83_2084) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2084;
      ov(63 downto 0) := iv;
      ptr_deref_2105_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2105_root_address_inst
    process(ptr_deref_2105_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2105_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2105_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2123_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2122;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2123_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2123_branch_req_0,
          ack0 => if_stmt_2123_branch_ack_0,
          ack1 => if_stmt_2123_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2174_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2173;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2174_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2174_branch_req_0,
          ack0 => if_stmt_2174_branch_ack_0,
          ack1 => if_stmt_2174_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1931_inst
    process(call7_1873) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1873, type_cast_1930_wire_constant, tmp_var);
      add45_1932 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1942_inst
    process(call9_1876) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1876, type_cast_1941_wire_constant, tmp_var);
      add58_1943 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2020_inst
    process(sub_1937, mul_2016) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1937, mul_2016, tmp_var);
      sub48_2021 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2030_inst
    process(sub61_1948, mul54_2026) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1948, mul54_2026, tmp_var);
      sub62_2031 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2134_inst
    process(input_dim2x_x1_1980) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1980, type_cast_2133_wire_constant, tmp_var);
      add98_2135 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2142_inst
    process(input_dim1x_x1_1987) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1987, type_cast_2141_wire_constant, tmp_var);
      inc_2143 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2156_inst
    process(inc110_2152, input_dim0x_x2_1994) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2152, input_dim0x_x2_1994, tmp_var);
      inc110x_xinput_dim0x_x2_2157 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2010_inst
    process(add_1910, tmp1_2006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1910, tmp1_2006, tmp_var);
      add_src_0x_x0_2011 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2116_inst
    process(conv90_2111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2111, type_cast_2115_wire_constant, tmp_var);
      add91_2117 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2205_inst
    process(indvar_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1973, type_cast_2204_wire_constant, tmp_var);
      indvarx_xnext_2206 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2052_inst
    process(mul76_2048, conv70_2039) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2048, conv70_2039, tmp_var);
      add77_2053 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2062_inst
    process(mul78_2058, conv65_2035) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2058, conv65_2035, tmp_var);
      add79_2063 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2095_inst
    process(shr85_2090) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2090, type_cast_2094_wire_constant, tmp_var);
      idxprom86_2096 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2147_inst
    process(inc_2143, call1_1864) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2143, call1_1864, tmp_var);
      cmp106_2148 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2172_inst
    process(conv112_2168, shr116132_1970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2168, shr116132_1970, tmp_var);
      cmp117_2173 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1925_inst
    process(call_1861) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1861, type_cast_1924_wire_constant, tmp_var);
      shr131_1926 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1969_inst
    process(conv115_1964) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1964, type_cast_1968_wire_constant, tmp_var);
      shr116132_1970 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2068_inst
    process(add_src_0x_x0_2011) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2011, type_cast_2067_wire_constant, tmp_var);
      shr81_2069 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2089_inst
    process(add79_2063) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2063, type_cast_2088_wire_constant, tmp_var);
      shr85_2090 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2015_inst
    process(input_dim0x_x2_1994, call13_1882) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1994, call13_1882, tmp_var);
      mul_2016 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2025_inst
    process(input_dim1x_x1_1987, call13_1882) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1987, call13_1882, tmp_var);
      mul54_2026 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2005_inst
    process(indvar_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1973, type_cast_2004_wire_constant, tmp_var);
      tmp1_2006 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2047_inst
    process(conv75_2043, conv73_1956) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2043, conv73_1956, tmp_var);
      mul76_2048 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2057_inst
    process(add77_2053, conv68_1952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2053, conv68_1952, tmp_var);
      mul78_2058 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1909_inst
    process(shl_1898, conv17_1905) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1898, conv17_1905, tmp_var);
      add_1910 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1897_inst
    process(conv_1892) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1892, type_cast_1896_wire_constant, tmp_var);
      shl_1898 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1936_inst
    process(add45_1932, call14_1885) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1932, call14_1885, tmp_var);
      sub_1937 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1947_inst
    process(add58_1943, call14_1885) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1943, call14_1885, tmp_var);
      sub61_1948 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2121_inst
    process(add91_2117, conv94_1960) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2117, conv94_1960, tmp_var);
      cmp_2122 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2078_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2077_scaled;
      array_obj_ref_2078_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2078_index_offset_req_0;
      array_obj_ref_2078_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2078_index_offset_req_1;
      array_obj_ref_2078_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2101_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2100_scaled;
      array_obj_ref_2101_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2101_index_offset_req_0;
      array_obj_ref_2101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2101_index_offset_req_1;
      array_obj_ref_2101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2083_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2083_load_0_req_0;
      ptr_deref_2083_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2083_load_0_req_1;
      ptr_deref_2083_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2083_word_address_0;
      ptr_deref_2083_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2105_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2105_store_0_req_0;
      ptr_deref_2105_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2105_store_0_req_1;
      ptr_deref_2105_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2105_word_address_0;
      data_in <= ptr_deref_2105_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1863_inst RPIPE_Block1_start_1860_inst RPIPE_Block1_start_1918_inst RPIPE_Block1_start_1915_inst RPIPE_Block1_start_1912_inst RPIPE_Block1_start_1900_inst RPIPE_Block1_start_1887_inst RPIPE_Block1_start_1884_inst RPIPE_Block1_start_1881_inst RPIPE_Block1_start_1878_inst RPIPE_Block1_start_1875_inst RPIPE_Block1_start_1872_inst RPIPE_Block1_start_1869_inst RPIPE_Block1_start_1866_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1863_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1860_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1918_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1915_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1912_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1900_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1887_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1884_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1881_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1878_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1875_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1872_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1869_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1866_inst_req_0;
      RPIPE_Block1_start_1863_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1860_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1918_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1915_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1912_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1900_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1887_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1884_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1881_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1878_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1875_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1872_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1869_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1866_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1863_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1860_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1918_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1915_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1912_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1900_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1887_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1884_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1881_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1878_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1875_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1872_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1869_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1866_inst_req_1;
      RPIPE_Block1_start_1863_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1860_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1918_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1915_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1912_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1900_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1887_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1884_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1881_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1878_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1875_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1872_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1869_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1866_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call1_1864 <= data_out(223 downto 208);
      call_1861 <= data_out(207 downto 192);
      call22_1919 <= data_out(191 downto 176);
      call20_1916 <= data_out(175 downto 160);
      call18_1913 <= data_out(159 downto 144);
      call16_1901 <= data_out(143 downto 128);
      call15_1888 <= data_out(127 downto 112);
      call14_1885 <= data_out(111 downto 96);
      call13_1882 <= data_out(95 downto 80);
      call11_1879 <= data_out(79 downto 64);
      call9_1876 <= data_out(63 downto 48);
      call7_1873 <= data_out(47 downto 32);
      call5_1870 <= data_out(31 downto 16);
      call3_1867 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2210_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2210_inst_req_0;
      WPIPE_Block1_done_2210_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2210_inst_req_1;
      WPIPE_Block1_done_2210_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2212_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5782_start: Boolean;
  signal convTransposeC_CP_5782_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2236_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2242_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2233_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2242_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2245_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2227_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2261_inst_req_1 : boolean;
  signal type_cast_2252_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2236_inst_req_1 : boolean;
  signal type_cast_2265_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2242_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2273_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2242_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2227_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2236_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2273_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2248_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2248_inst_ack_0 : boolean;
  signal type_cast_2252_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2233_inst_req_1 : boolean;
  signal type_cast_2265_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2261_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2230_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2233_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2248_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2233_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2239_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2279_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2230_inst_ack_1 : boolean;
  signal type_cast_2252_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2248_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2245_inst_req_0 : boolean;
  signal type_cast_2252_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2273_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2239_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2239_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2261_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2261_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2245_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2276_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2273_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2236_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2239_inst_ack_1 : boolean;
  signal type_cast_2265_inst_req_1 : boolean;
  signal type_cast_2265_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2227_inst_req_1 : boolean;
  signal type_cast_2312_inst_req_0 : boolean;
  signal type_cast_2312_inst_ack_0 : boolean;
  signal type_cast_2312_inst_req_1 : boolean;
  signal type_cast_2312_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2245_inst_ack_0 : boolean;
  signal type_cast_2320_inst_req_0 : boolean;
  signal type_cast_2320_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2279_inst_ack_1 : boolean;
  signal type_cast_2316_inst_req_1 : boolean;
  signal type_cast_2316_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2279_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2276_inst_ack_0 : boolean;
  signal type_cast_2316_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2276_inst_req_0 : boolean;
  signal type_cast_2316_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2279_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2230_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2230_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2227_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2276_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2221_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2221_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2221_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2221_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2224_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2224_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2224_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2224_inst_ack_1 : boolean;
  signal type_cast_2320_inst_req_1 : boolean;
  signal type_cast_2320_inst_ack_1 : boolean;
  signal type_cast_2324_inst_req_0 : boolean;
  signal type_cast_2324_inst_ack_0 : boolean;
  signal type_cast_2324_inst_req_1 : boolean;
  signal type_cast_2324_inst_ack_1 : boolean;
  signal type_cast_2406_inst_req_0 : boolean;
  signal type_cast_2406_inst_ack_0 : boolean;
  signal type_cast_2406_inst_req_1 : boolean;
  signal type_cast_2406_inst_ack_1 : boolean;
  signal type_cast_2410_inst_req_0 : boolean;
  signal type_cast_2410_inst_ack_0 : boolean;
  signal type_cast_2410_inst_req_1 : boolean;
  signal type_cast_2410_inst_ack_1 : boolean;
  signal type_cast_2414_inst_req_0 : boolean;
  signal type_cast_2414_inst_ack_0 : boolean;
  signal type_cast_2414_inst_req_1 : boolean;
  signal type_cast_2414_inst_ack_1 : boolean;
  signal type_cast_2444_inst_req_0 : boolean;
  signal type_cast_2444_inst_ack_0 : boolean;
  signal type_cast_2444_inst_req_1 : boolean;
  signal type_cast_2444_inst_ack_1 : boolean;
  signal array_obj_ref_2450_index_offset_req_0 : boolean;
  signal array_obj_ref_2450_index_offset_ack_0 : boolean;
  signal array_obj_ref_2450_index_offset_req_1 : boolean;
  signal array_obj_ref_2450_index_offset_ack_1 : boolean;
  signal addr_of_2451_final_reg_req_0 : boolean;
  signal addr_of_2451_final_reg_ack_0 : boolean;
  signal addr_of_2451_final_reg_req_1 : boolean;
  signal addr_of_2451_final_reg_ack_1 : boolean;
  signal ptr_deref_2455_load_0_req_0 : boolean;
  signal ptr_deref_2455_load_0_ack_0 : boolean;
  signal ptr_deref_2455_load_0_req_1 : boolean;
  signal ptr_deref_2455_load_0_ack_1 : boolean;
  signal array_obj_ref_2473_index_offset_req_0 : boolean;
  signal array_obj_ref_2473_index_offset_ack_0 : boolean;
  signal array_obj_ref_2473_index_offset_req_1 : boolean;
  signal array_obj_ref_2473_index_offset_ack_1 : boolean;
  signal addr_of_2474_final_reg_req_0 : boolean;
  signal addr_of_2474_final_reg_ack_0 : boolean;
  signal addr_of_2474_final_reg_req_1 : boolean;
  signal addr_of_2474_final_reg_ack_1 : boolean;
  signal ptr_deref_2477_store_0_req_0 : boolean;
  signal ptr_deref_2477_store_0_ack_0 : boolean;
  signal ptr_deref_2477_store_0_req_1 : boolean;
  signal ptr_deref_2477_store_0_ack_1 : boolean;
  signal type_cast_2482_inst_req_0 : boolean;
  signal type_cast_2482_inst_ack_0 : boolean;
  signal type_cast_2482_inst_req_1 : boolean;
  signal type_cast_2482_inst_ack_1 : boolean;
  signal if_stmt_2495_branch_req_0 : boolean;
  signal if_stmt_2495_branch_ack_1 : boolean;
  signal if_stmt_2495_branch_ack_0 : boolean;
  signal type_cast_2523_inst_req_0 : boolean;
  signal type_cast_2523_inst_ack_0 : boolean;
  signal type_cast_2523_inst_req_1 : boolean;
  signal type_cast_2523_inst_ack_1 : boolean;
  signal type_cast_2539_inst_req_0 : boolean;
  signal type_cast_2539_inst_ack_0 : boolean;
  signal type_cast_2539_inst_req_1 : boolean;
  signal type_cast_2539_inst_ack_1 : boolean;
  signal if_stmt_2546_branch_req_0 : boolean;
  signal if_stmt_2546_branch_ack_1 : boolean;
  signal if_stmt_2546_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2582_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2582_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2582_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2582_inst_ack_1 : boolean;
  signal phi_stmt_2345_req_0 : boolean;
  signal phi_stmt_2352_req_1 : boolean;
  signal phi_stmt_2359_req_1 : boolean;
  signal type_cast_2369_inst_req_0 : boolean;
  signal type_cast_2369_inst_ack_0 : boolean;
  signal type_cast_2369_inst_req_1 : boolean;
  signal type_cast_2369_inst_ack_1 : boolean;
  signal phi_stmt_2366_req_0 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal phi_stmt_2345_req_1 : boolean;
  signal type_cast_2355_inst_req_0 : boolean;
  signal type_cast_2355_inst_ack_0 : boolean;
  signal type_cast_2355_inst_req_1 : boolean;
  signal type_cast_2355_inst_ack_1 : boolean;
  signal phi_stmt_2352_req_0 : boolean;
  signal type_cast_2362_inst_req_0 : boolean;
  signal type_cast_2362_inst_ack_0 : boolean;
  signal type_cast_2362_inst_req_1 : boolean;
  signal type_cast_2362_inst_ack_1 : boolean;
  signal phi_stmt_2359_req_0 : boolean;
  signal type_cast_2371_inst_req_0 : boolean;
  signal type_cast_2371_inst_ack_0 : boolean;
  signal type_cast_2371_inst_req_1 : boolean;
  signal type_cast_2371_inst_ack_1 : boolean;
  signal phi_stmt_2366_req_1 : boolean;
  signal phi_stmt_2345_ack_0 : boolean;
  signal phi_stmt_2352_ack_0 : boolean;
  signal phi_stmt_2359_ack_0 : boolean;
  signal phi_stmt_2366_ack_0 : boolean;
  signal phi_stmt_2553_req_1 : boolean;
  signal type_cast_2565_inst_req_0 : boolean;
  signal type_cast_2565_inst_ack_0 : boolean;
  signal type_cast_2565_inst_req_1 : boolean;
  signal type_cast_2565_inst_ack_1 : boolean;
  signal phi_stmt_2560_req_1 : boolean;
  signal type_cast_2569_inst_req_0 : boolean;
  signal type_cast_2569_inst_ack_0 : boolean;
  signal type_cast_2569_inst_req_1 : boolean;
  signal type_cast_2569_inst_ack_1 : boolean;
  signal phi_stmt_2566_req_0 : boolean;
  signal type_cast_2556_inst_req_0 : boolean;
  signal type_cast_2556_inst_ack_0 : boolean;
  signal type_cast_2556_inst_req_1 : boolean;
  signal type_cast_2556_inst_ack_1 : boolean;
  signal phi_stmt_2553_req_0 : boolean;
  signal type_cast_2563_inst_req_0 : boolean;
  signal type_cast_2563_inst_ack_0 : boolean;
  signal type_cast_2563_inst_req_1 : boolean;
  signal type_cast_2563_inst_ack_1 : boolean;
  signal phi_stmt_2560_req_0 : boolean;
  signal type_cast_2571_inst_req_0 : boolean;
  signal type_cast_2571_inst_ack_0 : boolean;
  signal type_cast_2571_inst_req_1 : boolean;
  signal type_cast_2571_inst_ack_1 : boolean;
  signal phi_stmt_2566_req_1 : boolean;
  signal phi_stmt_2553_ack_0 : boolean;
  signal phi_stmt_2560_ack_0 : boolean;
  signal phi_stmt_2566_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5782_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5782_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5782_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5782_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5782: Block -- control-path 
    signal convTransposeC_CP_5782_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5782_elements(0) <= convTransposeC_CP_5782_start;
    convTransposeC_CP_5782_symbol <= convTransposeC_CP_5782_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2219/$entry
      -- CP-element group 0: 	 branch_block_stmt_2219/branch_block_stmt_2219__entry__
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280__entry__
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/$entry
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Sample/rr
      -- 
    cr_5975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(0), ack => type_cast_2252_inst_req_1); -- 
    cr_6003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(0), ack => type_cast_2265_inst_req_1); -- 
    rr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(0), ack => RPIPE_Block2_start_2221_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2219/merge_stmt_2552__exit__
      -- CP-element group 1: 	 branch_block_stmt_2219/assign_stmt_2578__entry__
      -- CP-element group 1: 	 branch_block_stmt_2219/assign_stmt_2578__exit__
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2219/assign_stmt_2578/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/assign_stmt_2578/$exit
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Update/cr
      -- 
    rr_6531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2351_inst_req_0); -- 
    cr_6536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2351_inst_req_1); -- 
    rr_6554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2355_inst_req_0); -- 
    cr_6559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2355_inst_req_1); -- 
    rr_6577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2362_inst_req_0); -- 
    cr_6582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2362_inst_req_1); -- 
    rr_6600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2371_inst_req_0); -- 
    cr_6605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(1), ack => type_cast_2371_inst_req_1); -- 
    convTransposeC_CP_5782_elements(1) <= convTransposeC_CP_5782_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Update/cr
      -- 
    ra_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2221_inst_ack_0, ack => convTransposeC_CP_5782_elements(2)); -- 
    cr_5835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(2), ack => RPIPE_Block2_start_2221_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2221_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Sample/rr
      -- 
    ca_5836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2221_inst_ack_1, ack => convTransposeC_CP_5782_elements(3)); -- 
    rr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(3), ack => RPIPE_Block2_start_2224_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Update/cr
      -- 
    ra_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2224_inst_ack_0, ack => convTransposeC_CP_5782_elements(4)); -- 
    cr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(4), ack => RPIPE_Block2_start_2224_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2224_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_sample_start_
      -- 
    ca_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2224_inst_ack_1, ack => convTransposeC_CP_5782_elements(5)); -- 
    rr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(5), ack => RPIPE_Block2_start_2227_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_update_start_
      -- 
    ra_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2227_inst_ack_0, ack => convTransposeC_CP_5782_elements(6)); -- 
    cr_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(6), ack => RPIPE_Block2_start_2227_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2227_update_completed_
      -- 
    ca_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2227_inst_ack_1, ack => convTransposeC_CP_5782_elements(7)); -- 
    rr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(7), ack => RPIPE_Block2_start_2230_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Sample/$exit
      -- 
    ra_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2230_inst_ack_0, ack => convTransposeC_CP_5782_elements(8)); -- 
    cr_5877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(8), ack => RPIPE_Block2_start_2230_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2230_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_sample_start_
      -- 
    ca_5878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2230_inst_ack_1, ack => convTransposeC_CP_5782_elements(9)); -- 
    rr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(9), ack => RPIPE_Block2_start_2233_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Update/cr
      -- 
    ra_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2233_inst_ack_0, ack => convTransposeC_CP_5782_elements(10)); -- 
    cr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(10), ack => RPIPE_Block2_start_2233_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2233_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Sample/rr
      -- 
    ca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2233_inst_ack_1, ack => convTransposeC_CP_5782_elements(11)); -- 
    rr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(11), ack => RPIPE_Block2_start_2236_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_sample_completed_
      -- 
    ra_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2236_inst_ack_0, ack => convTransposeC_CP_5782_elements(12)); -- 
    cr_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(12), ack => RPIPE_Block2_start_2236_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2236_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Sample/$entry
      -- 
    ca_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2236_inst_ack_1, ack => convTransposeC_CP_5782_elements(13)); -- 
    rr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(13), ack => RPIPE_Block2_start_2239_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Sample/$exit
      -- 
    ra_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2239_inst_ack_0, ack => convTransposeC_CP_5782_elements(14)); -- 
    cr_5919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(14), ack => RPIPE_Block2_start_2239_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2239_Update/$exit
      -- 
    ca_5920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2239_inst_ack_1, ack => convTransposeC_CP_5782_elements(15)); -- 
    rr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(15), ack => RPIPE_Block2_start_2242_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Sample/$exit
      -- 
    ra_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2242_inst_ack_0, ack => convTransposeC_CP_5782_elements(16)); -- 
    cr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(16), ack => RPIPE_Block2_start_2242_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2242_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_sample_start_
      -- 
    ca_5934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2242_inst_ack_1, ack => convTransposeC_CP_5782_elements(17)); -- 
    rr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(17), ack => RPIPE_Block2_start_2245_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Sample/ra
      -- 
    ra_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2245_inst_ack_0, ack => convTransposeC_CP_5782_elements(18)); -- 
    cr_5947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(18), ack => RPIPE_Block2_start_2245_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2245_Update/$exit
      -- 
    ca_5948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2245_inst_ack_1, ack => convTransposeC_CP_5782_elements(19)); -- 
    rr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(19), ack => RPIPE_Block2_start_2248_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Update/cr
      -- 
    ra_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2248_inst_ack_0, ack => convTransposeC_CP_5782_elements(20)); -- 
    cr_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(20), ack => RPIPE_Block2_start_2248_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2248_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Sample/$entry
      -- 
    ca_5962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2248_inst_ack_1, ack => convTransposeC_CP_5782_elements(21)); -- 
    rr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(21), ack => type_cast_2252_inst_req_0); -- 
    rr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(21), ack => RPIPE_Block2_start_2261_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Sample/$exit
      -- 
    ra_5971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_0, ack => convTransposeC_CP_5782_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2252_update_completed_
      -- 
    ca_5976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2252_inst_ack_1, ack => convTransposeC_CP_5782_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_sample_completed_
      -- 
    ra_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2261_inst_ack_0, ack => convTransposeC_CP_5782_elements(24)); -- 
    cr_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(24), ack => RPIPE_Block2_start_2261_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2261_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_sample_start_
      -- 
    ca_5990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2261_inst_ack_1, ack => convTransposeC_CP_5782_elements(25)); -- 
    rr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(25), ack => type_cast_2265_inst_req_0); -- 
    rr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(25), ack => RPIPE_Block2_start_2273_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_sample_completed_
      -- 
    ra_5999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2265_inst_ack_0, ack => convTransposeC_CP_5782_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/type_cast_2265_Update/ca
      -- 
    ca_6004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2265_inst_ack_1, ack => convTransposeC_CP_5782_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_sample_completed_
      -- 
    ra_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2273_inst_ack_0, ack => convTransposeC_CP_5782_elements(28)); -- 
    cr_6017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(28), ack => RPIPE_Block2_start_2273_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2273_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Sample/$entry
      -- 
    ca_6018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2273_inst_ack_1, ack => convTransposeC_CP_5782_elements(29)); -- 
    rr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(29), ack => RPIPE_Block2_start_2276_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_update_start_
      -- 
    ra_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2276_inst_ack_0, ack => convTransposeC_CP_5782_elements(30)); -- 
    cr_6031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(30), ack => RPIPE_Block2_start_2276_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2276_Update/ca
      -- 
    ca_6032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2276_inst_ack_1, ack => convTransposeC_CP_5782_elements(31)); -- 
    rr_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(31), ack => RPIPE_Block2_start_2279_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_sample_completed_
      -- 
    ra_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2279_inst_ack_0, ack => convTransposeC_CP_5782_elements(32)); -- 
    cr_6045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(32), ack => RPIPE_Block2_start_2279_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/RPIPE_Block2_start_2279_Update/$exit
      -- 
    ca_6046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2279_inst_ack_1, ack => convTransposeC_CP_5782_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280__exit__
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342__entry__
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2222_to_assign_stmt_2280/$exit
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Update/cr
      -- 
    rr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2312_inst_req_0); -- 
    cr_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2312_inst_req_1); -- 
    rr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2320_inst_req_0); -- 
    cr_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2316_inst_req_1); -- 
    rr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2316_inst_req_0); -- 
    cr_6090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2320_inst_req_1); -- 
    rr_6099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2324_inst_req_0); -- 
    cr_6104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(34), ack => type_cast_2324_inst_req_1); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(23) & convTransposeC_CP_5782_elements(27) & convTransposeC_CP_5782_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_sample_completed_
      -- 
    ra_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_0, ack => convTransposeC_CP_5782_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2312_Update/$exit
      -- 
    ca_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_1, ack => convTransposeC_CP_5782_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Sample/$exit
      -- 
    ra_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2316_inst_ack_0, ack => convTransposeC_CP_5782_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2316_Update/$exit
      -- 
    ca_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2316_inst_ack_1, ack => convTransposeC_CP_5782_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Sample/$exit
      -- 
    ra_6086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2320_inst_ack_0, ack => convTransposeC_CP_5782_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2320_Update/ca
      -- 
    ca_6091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2320_inst_ack_1, ack => convTransposeC_CP_5782_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Sample/ra
      -- 
    ra_6100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2324_inst_ack_0, ack => convTransposeC_CP_5782_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/type_cast_2324_Update/ca
      -- 
    ca_6105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2324_inst_ack_1, ack => convTransposeC_CP_5782_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342/$exit
      -- CP-element group 43: 	 branch_block_stmt_2219/assign_stmt_2287_to_assign_stmt_2342__exit__
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2345/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2352/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2359/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Update/cr
      -- 
    rr_6505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(43), ack => type_cast_2369_inst_req_0); -- 
    cr_6510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(43), ack => type_cast_2369_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(36) & convTransposeC_CP_5782_elements(38) & convTransposeC_CP_5782_elements(40) & convTransposeC_CP_5782_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Sample/ra
      -- 
    ra_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2406_inst_ack_0, ack => convTransposeC_CP_5782_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Update/ca
      -- 
    ca_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2406_inst_ack_1, ack => convTransposeC_CP_5782_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Sample/ra
      -- 
    ra_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2410_inst_ack_0, ack => convTransposeC_CP_5782_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Update/ca
      -- 
    ca_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2410_inst_ack_1, ack => convTransposeC_CP_5782_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Sample/ra
      -- 
    ra_6145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2414_inst_ack_0, ack => convTransposeC_CP_5782_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Update/ca
      -- 
    ca_6150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2414_inst_ack_1, ack => convTransposeC_CP_5782_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Sample/ra
      -- 
    ra_6159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2444_inst_ack_0, ack => convTransposeC_CP_5782_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Sample/req
      -- 
    ca_6164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2444_inst_ack_1, ack => convTransposeC_CP_5782_elements(51)); -- 
    req_6189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(51), ack => array_obj_ref_2450_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Sample/ack
      -- 
    ack_6190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2450_index_offset_ack_0, ack => convTransposeC_CP_5782_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_request/req
      -- 
    ack_6195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2450_index_offset_ack_1, ack => convTransposeC_CP_5782_elements(53)); -- 
    req_6204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(53), ack => addr_of_2451_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_request/ack
      -- 
    ack_6205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2451_final_reg_ack_0, ack => convTransposeC_CP_5782_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/word_access_start/word_0/rr
      -- 
    ack_6210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2451_final_reg_ack_1, ack => convTransposeC_CP_5782_elements(55)); -- 
    rr_6243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(55), ack => ptr_deref_2455_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Sample/word_access_start/word_0/ra
      -- 
    ra_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_0_ack_0, ack => convTransposeC_CP_5782_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/ptr_deref_2455_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/ptr_deref_2455_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/ptr_deref_2455_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/ptr_deref_2455_Merge/merge_ack
      -- 
    ca_6255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2455_load_0_ack_1, ack => convTransposeC_CP_5782_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Sample/req
      -- 
    req_6285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(58), ack => array_obj_ref_2473_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(45) & convTransposeC_CP_5782_elements(47) & convTransposeC_CP_5782_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Sample/ack
      -- 
    ack_6286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2473_index_offset_ack_0, ack => convTransposeC_CP_5782_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_request/req
      -- 
    ack_6291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2473_index_offset_ack_1, ack => convTransposeC_CP_5782_elements(60)); -- 
    req_6300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(60), ack => addr_of_2474_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_request/ack
      -- 
    ack_6301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2474_final_reg_ack_0, ack => convTransposeC_CP_5782_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_word_addrgen/root_register_ack
      -- 
    ack_6306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2474_final_reg_ack_1, ack => convTransposeC_CP_5782_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/ptr_deref_2477_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/ptr_deref_2477_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/ptr_deref_2477_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/ptr_deref_2477_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/word_access_start/word_0/rr
      -- 
    rr_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(63), ack => ptr_deref_2477_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(57) & convTransposeC_CP_5782_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Sample/word_access_start/word_0/ra
      -- 
    ra_6345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2477_store_0_ack_0, ack => convTransposeC_CP_5782_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/word_access_complete/word_0/ca
      -- 
    ca_6356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2477_store_0_ack_1, ack => convTransposeC_CP_5782_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Sample/ra
      -- 
    ra_6365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2482_inst_ack_0, ack => convTransposeC_CP_5782_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Update/ca
      -- 
    ca_6370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2482_inst_ack_1, ack => convTransposeC_CP_5782_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494__exit__
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495__entry__
      -- CP-element group 68: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/$exit
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2219/R_cmp_2496_place
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2219/if_stmt_2495_else_link/$entry
      -- 
    branch_req_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(68), ack => if_stmt_2495_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(52) & convTransposeC_CP_5782_elements(59) & convTransposeC_CP_5782_elements(65) & convTransposeC_CP_5782_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2219/merge_stmt_2501__exit__
      -- CP-element group 69: 	 branch_block_stmt_2219/assign_stmt_2507__entry__
      -- CP-element group 69: 	 branch_block_stmt_2219/assign_stmt_2507__exit__
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2219/if_stmt_2495_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2219/if_stmt_2495_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2219/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2219/assign_stmt_2507/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/assign_stmt_2507/$exit
      -- CP-element group 69: 	 branch_block_stmt_2219/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2219/merge_stmt_2501_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2219/merge_stmt_2501_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/merge_stmt_2501_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2219/merge_stmt_2501_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2495_branch_ack_1, ack => convTransposeC_CP_5782_elements(69)); -- 
    rr_6715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2556_inst_req_0); -- 
    cr_6720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2556_inst_req_1); -- 
    rr_6738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2563_inst_req_0); -- 
    cr_6743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2563_inst_req_1); -- 
    rr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2571_inst_req_0); -- 
    cr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(69), ack => type_cast_2571_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2219/merge_stmt_2509__exit__
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545__entry__
      -- CP-element group 70: 	 branch_block_stmt_2219/if_stmt_2495_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2219/if_stmt_2495_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2219/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/$entry
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2219/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2219/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2219/merge_stmt_2509_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2219/merge_stmt_2509_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2219/merge_stmt_2509_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2219/merge_stmt_2509_PhiAck/dummy
      -- 
    else_choice_transition_6387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2495_branch_ack_0, ack => convTransposeC_CP_5782_elements(70)); -- 
    rr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(70), ack => type_cast_2523_inst_req_0); -- 
    cr_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(70), ack => type_cast_2523_inst_req_1); -- 
    cr_6422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(70), ack => type_cast_2539_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Sample/ra
      -- 
    ra_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2523_inst_ack_0, ack => convTransposeC_CP_5782_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2523_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Sample/rr
      -- 
    ca_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2523_inst_ack_1, ack => convTransposeC_CP_5782_elements(72)); -- 
    rr_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(72), ack => type_cast_2539_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Sample/ra
      -- 
    ra_6418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2539_inst_ack_0, ack => convTransposeC_CP_5782_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545__exit__
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546__entry__
      -- CP-element group 74: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/$exit
      -- CP-element group 74: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2219/assign_stmt_2515_to_assign_stmt_2545/type_cast_2539_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2219/R_cmp122_2547_place
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2219/if_stmt_2546_else_link/$entry
      -- 
    ca_6423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2539_inst_ack_1, ack => convTransposeC_CP_5782_elements(74)); -- 
    branch_req_6431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(74), ack => if_stmt_2546_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2219/merge_stmt_2580__exit__
      -- CP-element group 75: 	 branch_block_stmt_2219/assign_stmt_2585__entry__
      -- CP-element group 75: 	 branch_block_stmt_2219/if_stmt_2546_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2219/if_stmt_2546_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2219/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2219/assign_stmt_2585/$entry
      -- CP-element group 75: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2219/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2219/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2219/merge_stmt_2580_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2219/merge_stmt_2580_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2219/merge_stmt_2580_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2219/merge_stmt_2580_PhiAck/dummy
      -- 
    if_choice_transition_6436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2546_branch_ack_1, ack => convTransposeC_CP_5782_elements(75)); -- 
    req_6456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(75), ack => WPIPE_Block2_done_2582_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2219/if_stmt_2546_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2219/if_stmt_2546_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2553/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2546_branch_ack_0, ack => convTransposeC_CP_5782_elements(76)); -- 
    rr_6666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2565_inst_req_0); -- 
    cr_6671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2565_inst_req_1); -- 
    rr_6689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2569_inst_req_0); -- 
    cr_6694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(76), ack => type_cast_2569_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Update/req
      -- 
    ack_6457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2582_inst_ack_0, ack => convTransposeC_CP_5782_elements(77)); -- 
    req_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(77), ack => WPIPE_Block2_done_2582_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2219/$exit
      -- CP-element group 78: 	 branch_block_stmt_2219/branch_block_stmt_2219__exit__
      -- CP-element group 78: 	 branch_block_stmt_2219/assign_stmt_2585__exit__
      -- CP-element group 78: 	 branch_block_stmt_2219/return__
      -- CP-element group 78: 	 branch_block_stmt_2219/merge_stmt_2587__exit__
      -- CP-element group 78: 	 branch_block_stmt_2219/assign_stmt_2585/$exit
      -- CP-element group 78: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2219/assign_stmt_2585/WPIPE_Block2_done_2582_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2219/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2219/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2219/merge_stmt_2587_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2219/merge_stmt_2587_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2219/merge_stmt_2587_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2219/merge_stmt_2587_PhiAck/dummy
      -- 
    ack_6462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2582_inst_ack_1, ack => convTransposeC_CP_5782_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2345/$exit
      -- CP-element group 79: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2349_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_req
      -- 
    phi_stmt_2345_req_6473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2345_req_6473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(79), ack => phi_stmt_2345_req_0); -- 
    -- Element group convTransposeC_CP_5782_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(43), ack => convTransposeC_CP_5782_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2352/$exit
      -- CP-element group 80: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2358_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_req
      -- 
    phi_stmt_2352_req_6481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2352_req_6481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(80), ack => phi_stmt_2352_req_1); -- 
    -- Element group convTransposeC_CP_5782_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(43), ack => convTransposeC_CP_5782_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2359/$exit
      -- CP-element group 81: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_req
      -- 
    phi_stmt_2359_req_6489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2359_req_6489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(81), ack => phi_stmt_2359_req_1); -- 
    -- Element group convTransposeC_CP_5782_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(43), ack => convTransposeC_CP_5782_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Sample/ra
      -- 
    ra_6506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2369_inst_ack_0, ack => convTransposeC_CP_5782_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/Update/ca
      -- 
    ca_6511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2369_inst_ack_1, ack => convTransposeC_CP_5782_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/$exit
      -- CP-element group 84: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/$exit
      -- CP-element group 84: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2369/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_req
      -- 
    phi_stmt_2366_req_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2366_req_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(84), ack => phi_stmt_2366_req_0); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(82) & convTransposeC_CP_5782_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2219/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(79) & convTransposeC_CP_5782_elements(80) & convTransposeC_CP_5782_elements(81) & convTransposeC_CP_5782_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Sample/ra
      -- 
    ra_6532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => convTransposeC_CP_5782_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/Update/ca
      -- 
    ca_6537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => convTransposeC_CP_5782_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/$exit
      -- CP-element group 88: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/$exit
      -- CP-element group 88: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_sources/type_cast_2351/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2345/phi_stmt_2345_req
      -- 
    phi_stmt_2345_req_6538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2345_req_6538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(88), ack => phi_stmt_2345_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(86) & convTransposeC_CP_5782_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Sample/ra
      -- 
    ra_6555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2355_inst_ack_0, ack => convTransposeC_CP_5782_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/Update/ca
      -- 
    ca_6560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2355_inst_ack_1, ack => convTransposeC_CP_5782_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/$exit
      -- CP-element group 91: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/$exit
      -- CP-element group 91: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_sources/type_cast_2355/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2352/phi_stmt_2352_req
      -- 
    phi_stmt_2352_req_6561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2352_req_6561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(91), ack => phi_stmt_2352_req_0); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(89) & convTransposeC_CP_5782_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Sample/ra
      -- 
    ra_6578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2362_inst_ack_0, ack => convTransposeC_CP_5782_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/Update/ca
      -- 
    ca_6583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2362_inst_ack_1, ack => convTransposeC_CP_5782_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/$exit
      -- CP-element group 94: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/$exit
      -- CP-element group 94: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2362/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_req
      -- 
    phi_stmt_2359_req_6584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2359_req_6584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(94), ack => phi_stmt_2359_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(92) & convTransposeC_CP_5782_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Sample/ra
      -- 
    ra_6601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_0, ack => convTransposeC_CP_5782_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/Update/ca
      -- 
    ca_6606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_1, ack => convTransposeC_CP_5782_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/$exit
      -- CP-element group 97: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/$exit
      -- CP-element group 97: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_sources/type_cast_2371/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2366/phi_stmt_2366_req
      -- 
    phi_stmt_2366_req_6607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2366_req_6607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(97), ack => phi_stmt_2366_req_1); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(95) & convTransposeC_CP_5782_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2219/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(88) & convTransposeC_CP_5782_elements(91) & convTransposeC_CP_5782_elements(94) & convTransposeC_CP_5782_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2219/merge_stmt_2344_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2219/merge_stmt_2344_PhiAck/$entry
      -- 
    convTransposeC_CP_5782_elements(99) <= OrReduce(convTransposeC_CP_5782_elements(85) & convTransposeC_CP_5782_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2219/merge_stmt_2344_PhiAck/phi_stmt_2345_ack
      -- 
    phi_stmt_2345_ack_6612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2345_ack_0, ack => convTransposeC_CP_5782_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2219/merge_stmt_2344_PhiAck/phi_stmt_2352_ack
      -- 
    phi_stmt_2352_ack_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2352_ack_0, ack => convTransposeC_CP_5782_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2219/merge_stmt_2344_PhiAck/phi_stmt_2359_ack
      -- 
    phi_stmt_2359_ack_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2359_ack_0, ack => convTransposeC_CP_5782_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2219/merge_stmt_2344_PhiAck/phi_stmt_2366_ack
      -- 
    phi_stmt_2366_ack_6615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2366_ack_0, ack => convTransposeC_CP_5782_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2219/merge_stmt_2344__exit__
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494__entry__
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2406_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2410_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2414_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2444_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2450_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2451_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2455_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/array_obj_ref_2473_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/addr_of_2474_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/ptr_deref_2477_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2219/assign_stmt_2378_to_assign_stmt_2494/type_cast_2482_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2219/merge_stmt_2344_PhiAck/$exit
      -- 
    rr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2406_inst_req_0); -- 
    cr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2406_inst_req_1); -- 
    rr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2410_inst_req_0); -- 
    cr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2410_inst_req_1); -- 
    rr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2414_inst_req_0); -- 
    cr_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2414_inst_req_1); -- 
    rr_6158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2444_inst_req_0); -- 
    cr_6163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2444_inst_req_1); -- 
    req_6194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => array_obj_ref_2450_index_offset_req_1); -- 
    req_6209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => addr_of_2451_final_reg_req_1); -- 
    cr_6254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => ptr_deref_2455_load_0_req_1); -- 
    req_6290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => array_obj_ref_2473_index_offset_req_1); -- 
    req_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => addr_of_2474_final_reg_req_1); -- 
    cr_6355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => ptr_deref_2477_store_0_req_1); -- 
    rr_6364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2482_inst_req_0); -- 
    cr_6369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(104), ack => type_cast_2482_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(100) & convTransposeC_CP_5782_elements(101) & convTransposeC_CP_5782_elements(102) & convTransposeC_CP_5782_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2553/$exit
      -- CP-element group 105: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_req
      -- 
    phi_stmt_2553_req_6650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2553_req_6650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(105), ack => phi_stmt_2553_req_1); -- 
    -- Element group convTransposeC_CP_5782_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5782_elements(76), ack => convTransposeC_CP_5782_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Sample/ra
      -- 
    ra_6667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_0, ack => convTransposeC_CP_5782_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/Update/ca
      -- 
    ca_6672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_1, ack => convTransposeC_CP_5782_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/$exit
      -- CP-element group 108: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/$exit
      -- CP-element group 108: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2565/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_req
      -- 
    phi_stmt_2560_req_6673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2560_req_6673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(108), ack => phi_stmt_2560_req_1); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(106) & convTransposeC_CP_5782_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Sample/ra
      -- 
    ra_6690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2569_inst_ack_0, ack => convTransposeC_CP_5782_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/Update/ca
      -- 
    ca_6695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2569_inst_ack_1, ack => convTransposeC_CP_5782_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/$exit
      -- CP-element group 111: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/$exit
      -- CP-element group 111: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2569/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_req
      -- 
    phi_stmt_2566_req_6696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2566_req_6696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(111), ack => phi_stmt_2566_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(109) & convTransposeC_CP_5782_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2219/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(105) & convTransposeC_CP_5782_elements(108) & convTransposeC_CP_5782_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Sample/ra
      -- 
    ra_6716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2556_inst_ack_0, ack => convTransposeC_CP_5782_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/Update/ca
      -- 
    ca_6721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2556_inst_ack_1, ack => convTransposeC_CP_5782_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/$exit
      -- CP-element group 115: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/$exit
      -- CP-element group 115: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2556/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2553/phi_stmt_2553_req
      -- 
    phi_stmt_2553_req_6722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2553_req_6722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(115), ack => phi_stmt_2553_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(113) & convTransposeC_CP_5782_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Sample/ra
      -- 
    ra_6739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2563_inst_ack_0, ack => convTransposeC_CP_5782_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/Update/ca
      -- 
    ca_6744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2563_inst_ack_1, ack => convTransposeC_CP_5782_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/$exit
      -- CP-element group 118: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/$exit
      -- CP-element group 118: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_sources/type_cast_2563/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2560/phi_stmt_2560_req
      -- 
    phi_stmt_2560_req_6745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2560_req_6745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(118), ack => phi_stmt_2560_req_0); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(116) & convTransposeC_CP_5782_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Sample/ra
      -- 
    ra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2571_inst_ack_0, ack => convTransposeC_CP_5782_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/Update/ca
      -- 
    ca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2571_inst_ack_1, ack => convTransposeC_CP_5782_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/$exit
      -- CP-element group 121: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/$exit
      -- CP-element group 121: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2571/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2566/phi_stmt_2566_req
      -- 
    phi_stmt_2566_req_6768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2566_req_6768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5782_elements(121), ack => phi_stmt_2566_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(119) & convTransposeC_CP_5782_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2219/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(115) & convTransposeC_CP_5782_elements(118) & convTransposeC_CP_5782_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2219/merge_stmt_2552_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2219/merge_stmt_2552_PhiAck/$entry
      -- 
    convTransposeC_CP_5782_elements(123) <= OrReduce(convTransposeC_CP_5782_elements(112) & convTransposeC_CP_5782_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2219/merge_stmt_2552_PhiAck/phi_stmt_2553_ack
      -- 
    phi_stmt_2553_ack_6773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2553_ack_0, ack => convTransposeC_CP_5782_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2219/merge_stmt_2552_PhiAck/phi_stmt_2560_ack
      -- 
    phi_stmt_2560_ack_6774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2560_ack_0, ack => convTransposeC_CP_5782_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2219/merge_stmt_2552_PhiAck/phi_stmt_2566_ack
      -- 
    phi_stmt_2566_ack_6775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2566_ack_0, ack => convTransposeC_CP_5782_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2219/merge_stmt_2552_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5782_elements(124) & convTransposeC_CP_5782_elements(125) & convTransposeC_CP_5782_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5782_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2472_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2472_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2449_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2449_scaled : std_logic_vector(13 downto 0);
    signal add121_2342 : std_logic_vector(31 downto 0);
    signal add45_2293 : std_logic_vector(15 downto 0);
    signal add58_2304 : std_logic_vector(15 downto 0);
    signal add77_2425 : std_logic_vector(63 downto 0);
    signal add79_2435 : std_logic_vector(63 downto 0);
    signal add91_2489 : std_logic_vector(31 downto 0);
    signal add98_2507 : std_logic_vector(15 downto 0);
    signal add_2271 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2383 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2450_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2450_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2450_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2450_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2450_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2450_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2473_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2473_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2473_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2473_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2473_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2473_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2452 : std_logic_vector(31 downto 0);
    signal arrayidx87_2475 : std_logic_vector(31 downto 0);
    signal call11_2240 : std_logic_vector(15 downto 0);
    signal call13_2243 : std_logic_vector(15 downto 0);
    signal call14_2246 : std_logic_vector(15 downto 0);
    signal call15_2249 : std_logic_vector(15 downto 0);
    signal call16_2262 : std_logic_vector(15 downto 0);
    signal call18_2274 : std_logic_vector(15 downto 0);
    signal call1_2225 : std_logic_vector(15 downto 0);
    signal call20_2277 : std_logic_vector(15 downto 0);
    signal call22_2280 : std_logic_vector(15 downto 0);
    signal call3_2228 : std_logic_vector(15 downto 0);
    signal call5_2231 : std_logic_vector(15 downto 0);
    signal call7_2234 : std_logic_vector(15 downto 0);
    signal call9_2237 : std_logic_vector(15 downto 0);
    signal call_2222 : std_logic_vector(15 downto 0);
    signal cmp106_2520 : std_logic_vector(0 downto 0);
    signal cmp122_2545 : std_logic_vector(0 downto 0);
    signal cmp_2494 : std_logic_vector(0 downto 0);
    signal conv112_2540 : std_logic_vector(31 downto 0);
    signal conv115_2325 : std_logic_vector(31 downto 0);
    signal conv17_2266 : std_logic_vector(31 downto 0);
    signal conv65_2407 : std_logic_vector(63 downto 0);
    signal conv68_2313 : std_logic_vector(63 downto 0);
    signal conv70_2411 : std_logic_vector(63 downto 0);
    signal conv73_2317 : std_logic_vector(63 downto 0);
    signal conv75_2415 : std_logic_vector(63 downto 0);
    signal conv90_2483 : std_logic_vector(31 downto 0);
    signal conv94_2321 : std_logic_vector(31 downto 0);
    signal conv_2253 : std_logic_vector(31 downto 0);
    signal idxprom86_2468 : std_logic_vector(63 downto 0);
    signal idxprom_2445 : std_logic_vector(63 downto 0);
    signal inc110_2524 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2529 : std_logic_vector(15 downto 0);
    signal inc_2515 : std_logic_vector(15 downto 0);
    signal indvar_2345 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2578 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2566 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2366 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2560 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2359 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2536 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2553 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2352 : std_logic_vector(15 downto 0);
    signal mul54_2398 : std_logic_vector(15 downto 0);
    signal mul76_2420 : std_logic_vector(63 downto 0);
    signal mul78_2430 : std_logic_vector(63 downto 0);
    signal mul_2388 : std_logic_vector(15 downto 0);
    signal ptr_deref_2455_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2455_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2455_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2455_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2455_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2477_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2477_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2477_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2477_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2477_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2477_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2259 : std_logic_vector(31 downto 0);
    signal shr116137_2331 : std_logic_vector(31 downto 0);
    signal shr120138_2337 : std_logic_vector(31 downto 0);
    signal shr136_2287 : std_logic_vector(15 downto 0);
    signal shr81_2441 : std_logic_vector(31 downto 0);
    signal shr85_2462 : std_logic_vector(63 downto 0);
    signal sub48_2393 : std_logic_vector(15 downto 0);
    signal sub61_2309 : std_logic_vector(15 downto 0);
    signal sub62_2403 : std_logic_vector(15 downto 0);
    signal sub_2298 : std_logic_vector(15 downto 0);
    signal tmp1_2378 : std_logic_vector(31 downto 0);
    signal tmp83_2456 : std_logic_vector(63 downto 0);
    signal type_cast_2257_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2285_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2291_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2302_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2329_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2335_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2349_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2351_wire : std_logic_vector(31 downto 0);
    signal type_cast_2355_wire : std_logic_vector(15 downto 0);
    signal type_cast_2358_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2362_wire : std_logic_vector(15 downto 0);
    signal type_cast_2365_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2369_wire : std_logic_vector(15 downto 0);
    signal type_cast_2371_wire : std_logic_vector(15 downto 0);
    signal type_cast_2376_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2439_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2460_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2466_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2487_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2505_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2513_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2533_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2556_wire : std_logic_vector(15 downto 0);
    signal type_cast_2559_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2563_wire : std_logic_vector(15 downto 0);
    signal type_cast_2565_wire : std_logic_vector(15 downto 0);
    signal type_cast_2569_wire : std_logic_vector(15 downto 0);
    signal type_cast_2571_wire : std_logic_vector(15 downto 0);
    signal type_cast_2576_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2584_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2450_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2450_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2450_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2450_resized_base_address <= "00000000000000";
    array_obj_ref_2473_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2473_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2473_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2473_resized_base_address <= "00000000000000";
    ptr_deref_2455_word_offset_0 <= "00000000000000";
    ptr_deref_2477_word_offset_0 <= "00000000000000";
    type_cast_2257_wire_constant <= "00000000000000000000000000010000";
    type_cast_2285_wire_constant <= "0000000000000001";
    type_cast_2291_wire_constant <= "1111111111111111";
    type_cast_2302_wire_constant <= "1111111111111111";
    type_cast_2329_wire_constant <= "00000000000000000000000000000010";
    type_cast_2335_wire_constant <= "00000000000000000000000000000001";
    type_cast_2349_wire_constant <= "00000000000000000000000000000000";
    type_cast_2358_wire_constant <= "0000000000000000";
    type_cast_2365_wire_constant <= "0000000000000000";
    type_cast_2376_wire_constant <= "00000000000000000000000000000100";
    type_cast_2439_wire_constant <= "00000000000000000000000000000010";
    type_cast_2460_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2466_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2487_wire_constant <= "00000000000000000000000000000100";
    type_cast_2505_wire_constant <= "0000000000000100";
    type_cast_2513_wire_constant <= "0000000000000001";
    type_cast_2533_wire_constant <= "0000000000000000";
    type_cast_2559_wire_constant <= "0000000000000000";
    type_cast_2576_wire_constant <= "00000000000000000000000000000001";
    type_cast_2584_wire_constant <= "0000000000000001";
    phi_stmt_2345: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2349_wire_constant & type_cast_2351_wire;
      req <= phi_stmt_2345_req_0 & phi_stmt_2345_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2345",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2345_ack_0,
          idata => idata,
          odata => indvar_2345,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2345
    phi_stmt_2352: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2355_wire & type_cast_2358_wire_constant;
      req <= phi_stmt_2352_req_0 & phi_stmt_2352_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2352",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2352_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2352
    phi_stmt_2359: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2362_wire & type_cast_2365_wire_constant;
      req <= phi_stmt_2359_req_0 & phi_stmt_2359_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2359",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2359_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2359,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2359
    phi_stmt_2366: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2369_wire & type_cast_2371_wire;
      req <= phi_stmt_2366_req_0 & phi_stmt_2366_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2366",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2366_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2366,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2366
    phi_stmt_2553: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2556_wire & type_cast_2559_wire_constant;
      req <= phi_stmt_2553_req_0 & phi_stmt_2553_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2553",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2553_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2553,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2553
    phi_stmt_2560: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2563_wire & type_cast_2565_wire;
      req <= phi_stmt_2560_req_0 & phi_stmt_2560_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2560",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2560_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2560,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2560
    phi_stmt_2566: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2569_wire & type_cast_2571_wire;
      req <= phi_stmt_2566_req_0 & phi_stmt_2566_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2566",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2566_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2566,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2566
    -- flow-through select operator MUX_2535_inst
    input_dim1x_x2_2536 <= type_cast_2533_wire_constant when (cmp106_2520(0) /=  '0') else inc_2515;
    addr_of_2451_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2451_final_reg_req_0;
      addr_of_2451_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2451_final_reg_req_1;
      addr_of_2451_final_reg_ack_1<= rack(0);
      addr_of_2451_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2451_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2450_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2452,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2474_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2474_final_reg_req_0;
      addr_of_2474_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2474_final_reg_req_1;
      addr_of_2474_final_reg_ack_1<= rack(0);
      addr_of_2474_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2474_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2473_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2252_inst_req_0;
      type_cast_2252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2252_inst_req_1;
      type_cast_2252_inst_ack_1<= rack(0);
      type_cast_2252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2249,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2265_inst_req_0;
      type_cast_2265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2265_inst_req_1;
      type_cast_2265_inst_ack_1<= rack(0);
      type_cast_2265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2312_inst_req_0;
      type_cast_2312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2312_inst_req_1;
      type_cast_2312_inst_ack_1<= rack(0);
      type_cast_2312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2316_inst_req_0;
      type_cast_2316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2316_inst_req_1;
      type_cast_2316_inst_ack_1<= rack(0);
      type_cast_2316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2320_inst_req_0;
      type_cast_2320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2320_inst_req_1;
      type_cast_2320_inst_ack_1<= rack(0);
      type_cast_2320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2324_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2324_inst_req_0;
      type_cast_2324_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2324_inst_req_1;
      type_cast_2324_inst_ack_1<= rack(0);
      type_cast_2324_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2324_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2578,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2351_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2355_inst_req_0;
      type_cast_2355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2355_inst_req_1;
      type_cast_2355_inst_ack_1<= rack(0);
      type_cast_2355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2355_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2362_inst_req_0;
      type_cast_2362_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2362_inst_req_1;
      type_cast_2362_inst_ack_1<= rack(0);
      type_cast_2362_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2362_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2560,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2362_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2369_inst_req_0;
      type_cast_2369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2369_inst_req_1;
      type_cast_2369_inst_ack_1<= rack(0);
      type_cast_2369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2369_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2369_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2371_inst_req_0;
      type_cast_2371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2371_inst_req_1;
      type_cast_2371_inst_ack_1<= rack(0);
      type_cast_2371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2371_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2406_inst_req_0;
      type_cast_2406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2406_inst_req_1;
      type_cast_2406_inst_ack_1<= rack(0);
      type_cast_2406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2410_inst_req_0;
      type_cast_2410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2410_inst_req_1;
      type_cast_2410_inst_ack_1<= rack(0);
      type_cast_2410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2414_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2414_inst_req_0;
      type_cast_2414_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2414_inst_req_1;
      type_cast_2414_inst_ack_1<= rack(0);
      type_cast_2414_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2414_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2415,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2444_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2444_inst_req_0;
      type_cast_2444_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2444_inst_req_1;
      type_cast_2444_inst_ack_1<= rack(0);
      type_cast_2444_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2444_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2445,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2482_inst_req_0;
      type_cast_2482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2482_inst_req_1;
      type_cast_2482_inst_ack_1<= rack(0);
      type_cast_2482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2523_inst_req_0;
      type_cast_2523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2523_inst_req_1;
      type_cast_2523_inst_ack_1<= rack(0);
      type_cast_2523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2539_inst_req_0;
      type_cast_2539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2539_inst_req_1;
      type_cast_2539_inst_ack_1<= rack(0);
      type_cast_2539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2556_inst_req_0;
      type_cast_2556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2556_inst_req_1;
      type_cast_2556_inst_ack_1<= rack(0);
      type_cast_2556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2556_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2563_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2563_inst_req_0;
      type_cast_2563_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2563_inst_req_1;
      type_cast_2563_inst_ack_1<= rack(0);
      type_cast_2563_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2563_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2359,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2563_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2565_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2565_inst_req_0;
      type_cast_2565_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2565_inst_req_1;
      type_cast_2565_inst_ack_1<= rack(0);
      type_cast_2565_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2565_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2565_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2569_inst_req_0;
      type_cast_2569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2569_inst_req_1;
      type_cast_2569_inst_ack_1<= rack(0);
      type_cast_2569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2569_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2571_inst_req_0;
      type_cast_2571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2571_inst_req_1;
      type_cast_2571_inst_ack_1<= rack(0);
      type_cast_2571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2571_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2450_index_1_rename
    process(R_idxprom_2449_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2449_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2449_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2450_index_1_resize
    process(idxprom_2445) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2445;
      ov := iv(13 downto 0);
      R_idxprom_2449_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2450_root_address_inst
    process(array_obj_ref_2450_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2450_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2450_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2473_index_1_rename
    process(R_idxprom86_2472_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2472_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2472_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2473_index_1_resize
    process(idxprom86_2468) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2468;
      ov := iv(13 downto 0);
      R_idxprom86_2472_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2473_root_address_inst
    process(array_obj_ref_2473_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2473_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2473_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2455_addr_0
    process(ptr_deref_2455_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2455_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2455_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2455_base_resize
    process(arrayidx82_2452) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2452;
      ov := iv(13 downto 0);
      ptr_deref_2455_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2455_gather_scatter
    process(ptr_deref_2455_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2455_data_0;
      ov(63 downto 0) := iv;
      tmp83_2456 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2455_root_address_inst
    process(ptr_deref_2455_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2455_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2455_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2477_addr_0
    process(ptr_deref_2477_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2477_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2477_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2477_base_resize
    process(arrayidx87_2475) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2475;
      ov := iv(13 downto 0);
      ptr_deref_2477_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2477_gather_scatter
    process(tmp83_2456) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2456;
      ov(63 downto 0) := iv;
      ptr_deref_2477_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2477_root_address_inst
    process(ptr_deref_2477_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2477_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2477_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2495_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2494;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2495_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2495_branch_req_0,
          ack0 => if_stmt_2495_branch_ack_0,
          ack1 => if_stmt_2495_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2546_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2545;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2546_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2546_branch_req_0,
          ack0 => if_stmt_2546_branch_ack_0,
          ack1 => if_stmt_2546_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2292_inst
    process(call7_2234) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2234, type_cast_2291_wire_constant, tmp_var);
      add45_2293 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2303_inst
    process(call9_2237) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2237, type_cast_2302_wire_constant, tmp_var);
      add58_2304 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2392_inst
    process(sub_2298, mul_2388) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2298, mul_2388, tmp_var);
      sub48_2393 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2402_inst
    process(sub61_2309, mul54_2398) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2309, mul54_2398, tmp_var);
      sub62_2403 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2506_inst
    process(input_dim2x_x1_2352) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2352, type_cast_2505_wire_constant, tmp_var);
      add98_2507 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2514_inst
    process(input_dim1x_x1_2359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2359, type_cast_2513_wire_constant, tmp_var);
      inc_2515 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2528_inst
    process(inc110_2524, input_dim0x_x2_2366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2524, input_dim0x_x2_2366, tmp_var);
      inc110x_xinput_dim0x_x2_2529 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2341_inst
    process(shr116137_2331, shr120138_2337) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2331, shr120138_2337, tmp_var);
      add121_2342 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2382_inst
    process(add_2271, tmp1_2378) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2271, tmp1_2378, tmp_var);
      add_src_0x_x0_2383 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2488_inst
    process(conv90_2483) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2483, type_cast_2487_wire_constant, tmp_var);
      add91_2489 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2577_inst
    process(indvar_2345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2345, type_cast_2576_wire_constant, tmp_var);
      indvarx_xnext_2578 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2424_inst
    process(mul76_2420, conv70_2411) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2420, conv70_2411, tmp_var);
      add77_2425 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2434_inst
    process(mul78_2430, conv65_2407) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2430, conv65_2407, tmp_var);
      add79_2435 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2467_inst
    process(shr85_2462) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2462, type_cast_2466_wire_constant, tmp_var);
      idxprom86_2468 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2519_inst
    process(inc_2515, call1_2225) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2515, call1_2225, tmp_var);
      cmp106_2520 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2544_inst
    process(conv112_2540, add121_2342) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2540, add121_2342, tmp_var);
      cmp122_2545 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2286_inst
    process(call_2222) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2222, type_cast_2285_wire_constant, tmp_var);
      shr136_2287 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2330_inst
    process(conv115_2325) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2325, type_cast_2329_wire_constant, tmp_var);
      shr116137_2331 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2336_inst
    process(conv115_2325) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2325, type_cast_2335_wire_constant, tmp_var);
      shr120138_2337 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2440_inst
    process(add_src_0x_x0_2383) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2383, type_cast_2439_wire_constant, tmp_var);
      shr81_2441 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2461_inst
    process(add79_2435) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2435, type_cast_2460_wire_constant, tmp_var);
      shr85_2462 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2387_inst
    process(input_dim0x_x2_2366, call13_2243) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2366, call13_2243, tmp_var);
      mul_2388 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2397_inst
    process(input_dim1x_x1_2359, call13_2243) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2359, call13_2243, tmp_var);
      mul54_2398 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2377_inst
    process(indvar_2345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2345, type_cast_2376_wire_constant, tmp_var);
      tmp1_2378 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2419_inst
    process(conv75_2415, conv73_2317) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2415, conv73_2317, tmp_var);
      mul76_2420 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2429_inst
    process(add77_2425, conv68_2313) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2425, conv68_2313, tmp_var);
      mul78_2430 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2270_inst
    process(shl_2259, conv17_2266) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2259, conv17_2266, tmp_var);
      add_2271 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2258_inst
    process(conv_2253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2253, type_cast_2257_wire_constant, tmp_var);
      shl_2259 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2297_inst
    process(add45_2293, call14_2246) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2293, call14_2246, tmp_var);
      sub_2298 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2308_inst
    process(add58_2304, call14_2246) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2304, call14_2246, tmp_var);
      sub61_2309 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2493_inst
    process(add91_2489, conv94_2321) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2489, conv94_2321, tmp_var);
      cmp_2494 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2450_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2449_scaled;
      array_obj_ref_2450_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2450_index_offset_req_0;
      array_obj_ref_2450_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2450_index_offset_req_1;
      array_obj_ref_2450_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2473_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2472_scaled;
      array_obj_ref_2473_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2473_index_offset_req_0;
      array_obj_ref_2473_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2473_index_offset_req_1;
      array_obj_ref_2473_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2455_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2455_load_0_req_0;
      ptr_deref_2455_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2455_load_0_req_1;
      ptr_deref_2455_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2455_word_address_0;
      ptr_deref_2455_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2477_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2477_store_0_req_0;
      ptr_deref_2477_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2477_store_0_req_1;
      ptr_deref_2477_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2477_word_address_0;
      data_in <= ptr_deref_2477_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2245_inst RPIPE_Block2_start_2248_inst RPIPE_Block2_start_2261_inst RPIPE_Block2_start_2273_inst RPIPE_Block2_start_2276_inst RPIPE_Block2_start_2279_inst RPIPE_Block2_start_2242_inst RPIPE_Block2_start_2239_inst RPIPE_Block2_start_2236_inst RPIPE_Block2_start_2233_inst RPIPE_Block2_start_2230_inst RPIPE_Block2_start_2227_inst RPIPE_Block2_start_2224_inst RPIPE_Block2_start_2221_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2245_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2248_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2261_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2273_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2276_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2279_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2242_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2239_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2236_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2233_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2230_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2227_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2224_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2221_inst_req_0;
      RPIPE_Block2_start_2245_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2248_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2261_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2273_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2276_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2279_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2242_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2239_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2236_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2233_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2230_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2227_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2224_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2221_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2245_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2248_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2261_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2273_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2276_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2279_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2242_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2239_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2236_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2233_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2230_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2227_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2224_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2221_inst_req_1;
      RPIPE_Block2_start_2245_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2248_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2261_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2273_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2276_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2279_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2242_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2239_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2236_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2233_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2230_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2227_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2224_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2221_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call14_2246 <= data_out(223 downto 208);
      call15_2249 <= data_out(207 downto 192);
      call16_2262 <= data_out(191 downto 176);
      call18_2274 <= data_out(175 downto 160);
      call20_2277 <= data_out(159 downto 144);
      call22_2280 <= data_out(143 downto 128);
      call13_2243 <= data_out(127 downto 112);
      call11_2240 <= data_out(111 downto 96);
      call9_2237 <= data_out(95 downto 80);
      call7_2234 <= data_out(79 downto 64);
      call5_2231 <= data_out(63 downto 48);
      call3_2228 <= data_out(47 downto 32);
      call1_2225 <= data_out(31 downto 16);
      call_2222 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2582_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2582_inst_req_0;
      WPIPE_Block2_done_2582_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2582_inst_req_1;
      WPIPE_Block2_done_2582_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2584_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6792_start: Boolean;
  signal convTransposeD_CP_6792_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2593_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2593_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2645_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2614_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2617_inst_ack_0 : boolean;
  signal type_cast_2699_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2602_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2648_inst_ack_0 : boolean;
  signal type_cast_2695_inst_req_1 : boolean;
  signal type_cast_2695_inst_req_0 : boolean;
  signal type_cast_2768_inst_req_0 : boolean;
  signal type_cast_2768_inst_ack_0 : boolean;
  signal type_cast_2637_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2611_inst_req_1 : boolean;
  signal type_cast_2695_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2611_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2633_inst_ack_1 : boolean;
  signal type_cast_2695_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2620_inst_ack_1 : boolean;
  signal type_cast_2806_inst_req_1 : boolean;
  signal type_cast_2806_inst_ack_1 : boolean;
  signal type_cast_2768_inst_req_1 : boolean;
  signal type_cast_2768_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2605_inst_ack_1 : boolean;
  signal type_cast_2699_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2593_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2593_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2614_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2648_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2599_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2617_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2617_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2605_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2633_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2648_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2602_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2645_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2596_inst_req_1 : boolean;
  signal type_cast_2703_inst_req_0 : boolean;
  signal type_cast_2703_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2608_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2633_inst_req_0 : boolean;
  signal type_cast_2624_inst_req_1 : boolean;
  signal type_cast_2624_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2645_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2645_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2651_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2596_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2614_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2614_inst_ack_1 : boolean;
  signal type_cast_2624_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2651_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2648_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2633_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2617_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2596_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2596_inst_ack_0 : boolean;
  signal type_cast_2624_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2651_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2651_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2605_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2602_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2605_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2602_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2611_inst_ack_0 : boolean;
  signal type_cast_2703_inst_req_1 : boolean;
  signal type_cast_2703_inst_ack_1 : boolean;
  signal type_cast_2699_inst_ack_1 : boolean;
  signal type_cast_2699_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2611_inst_req_0 : boolean;
  signal type_cast_2776_inst_ack_1 : boolean;
  signal type_cast_2637_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2620_inst_req_1 : boolean;
  signal type_cast_2772_inst_ack_1 : boolean;
  signal type_cast_2637_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2620_inst_ack_0 : boolean;
  signal array_obj_ref_2812_index_offset_req_1 : boolean;
  signal array_obj_ref_2812_index_offset_ack_1 : boolean;
  signal type_cast_2776_inst_req_1 : boolean;
  signal type_cast_2637_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2620_inst_req_0 : boolean;
  signal addr_of_2813_final_reg_req_1 : boolean;
  signal addr_of_2813_final_reg_ack_1 : boolean;
  signal RPIPE_Block3_start_2608_inst_ack_1 : boolean;
  signal array_obj_ref_2812_index_offset_req_0 : boolean;
  signal array_obj_ref_2812_index_offset_ack_0 : boolean;
  signal RPIPE_Block3_start_2608_inst_req_1 : boolean;
  signal addr_of_2813_final_reg_req_0 : boolean;
  signal addr_of_2813_final_reg_ack_0 : boolean;
  signal type_cast_2806_inst_req_0 : boolean;
  signal type_cast_2806_inst_ack_0 : boolean;
  signal type_cast_2772_inst_req_0 : boolean;
  signal type_cast_2772_inst_ack_0 : boolean;
  signal type_cast_2776_inst_req_0 : boolean;
  signal type_cast_2776_inst_ack_0 : boolean;
  signal type_cast_2772_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2608_inst_ack_0 : boolean;
  signal ptr_deref_2817_load_0_req_0 : boolean;
  signal ptr_deref_2817_load_0_ack_0 : boolean;
  signal ptr_deref_2817_load_0_req_1 : boolean;
  signal ptr_deref_2817_load_0_ack_1 : boolean;
  signal array_obj_ref_2835_index_offset_req_0 : boolean;
  signal array_obj_ref_2835_index_offset_ack_0 : boolean;
  signal array_obj_ref_2835_index_offset_req_1 : boolean;
  signal array_obj_ref_2835_index_offset_ack_1 : boolean;
  signal addr_of_2836_final_reg_req_0 : boolean;
  signal addr_of_2836_final_reg_ack_0 : boolean;
  signal addr_of_2836_final_reg_req_1 : boolean;
  signal addr_of_2836_final_reg_ack_1 : boolean;
  signal ptr_deref_2839_store_0_req_0 : boolean;
  signal ptr_deref_2839_store_0_ack_0 : boolean;
  signal ptr_deref_2839_store_0_req_1 : boolean;
  signal ptr_deref_2839_store_0_ack_1 : boolean;
  signal type_cast_2844_inst_req_0 : boolean;
  signal type_cast_2844_inst_ack_0 : boolean;
  signal type_cast_2844_inst_req_1 : boolean;
  signal type_cast_2844_inst_ack_1 : boolean;
  signal if_stmt_2857_branch_req_0 : boolean;
  signal if_stmt_2857_branch_ack_1 : boolean;
  signal if_stmt_2857_branch_ack_0 : boolean;
  signal type_cast_2885_inst_req_0 : boolean;
  signal type_cast_2885_inst_ack_0 : boolean;
  signal type_cast_2885_inst_req_1 : boolean;
  signal type_cast_2885_inst_ack_1 : boolean;
  signal if_stmt_2904_branch_req_0 : boolean;
  signal if_stmt_2904_branch_ack_1 : boolean;
  signal if_stmt_2904_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2940_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2940_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2940_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2940_inst_ack_1 : boolean;
  signal phi_stmt_2707_req_0 : boolean;
  signal phi_stmt_2714_req_0 : boolean;
  signal phi_stmt_2721_req_0 : boolean;
  signal type_cast_2731_inst_req_0 : boolean;
  signal type_cast_2731_inst_ack_0 : boolean;
  signal type_cast_2731_inst_req_1 : boolean;
  signal type_cast_2731_inst_ack_1 : boolean;
  signal phi_stmt_2728_req_0 : boolean;
  signal type_cast_2713_inst_req_0 : boolean;
  signal type_cast_2713_inst_ack_0 : boolean;
  signal type_cast_2713_inst_req_1 : boolean;
  signal type_cast_2713_inst_ack_1 : boolean;
  signal phi_stmt_2707_req_1 : boolean;
  signal type_cast_2720_inst_req_0 : boolean;
  signal type_cast_2720_inst_ack_0 : boolean;
  signal type_cast_2720_inst_req_1 : boolean;
  signal type_cast_2720_inst_ack_1 : boolean;
  signal phi_stmt_2714_req_1 : boolean;
  signal type_cast_2727_inst_req_0 : boolean;
  signal type_cast_2727_inst_ack_0 : boolean;
  signal type_cast_2727_inst_req_1 : boolean;
  signal type_cast_2727_inst_ack_1 : boolean;
  signal phi_stmt_2721_req_1 : boolean;
  signal type_cast_2733_inst_req_0 : boolean;
  signal type_cast_2733_inst_ack_0 : boolean;
  signal type_cast_2733_inst_req_1 : boolean;
  signal type_cast_2733_inst_ack_1 : boolean;
  signal phi_stmt_2728_req_1 : boolean;
  signal phi_stmt_2707_ack_0 : boolean;
  signal phi_stmt_2714_ack_0 : boolean;
  signal phi_stmt_2721_ack_0 : boolean;
  signal phi_stmt_2728_ack_0 : boolean;
  signal phi_stmt_2911_req_1 : boolean;
  signal type_cast_2923_inst_req_0 : boolean;
  signal type_cast_2923_inst_ack_0 : boolean;
  signal type_cast_2923_inst_req_1 : boolean;
  signal type_cast_2923_inst_ack_1 : boolean;
  signal phi_stmt_2918_req_1 : boolean;
  signal type_cast_2929_inst_req_0 : boolean;
  signal type_cast_2929_inst_ack_0 : boolean;
  signal type_cast_2929_inst_req_1 : boolean;
  signal type_cast_2929_inst_ack_1 : boolean;
  signal phi_stmt_2924_req_1 : boolean;
  signal type_cast_2914_inst_req_0 : boolean;
  signal type_cast_2914_inst_ack_0 : boolean;
  signal type_cast_2914_inst_req_1 : boolean;
  signal type_cast_2914_inst_ack_1 : boolean;
  signal phi_stmt_2911_req_0 : boolean;
  signal type_cast_2921_inst_req_0 : boolean;
  signal type_cast_2921_inst_ack_0 : boolean;
  signal type_cast_2921_inst_req_1 : boolean;
  signal type_cast_2921_inst_ack_1 : boolean;
  signal phi_stmt_2918_req_0 : boolean;
  signal type_cast_2927_inst_req_0 : boolean;
  signal type_cast_2927_inst_ack_0 : boolean;
  signal type_cast_2927_inst_req_1 : boolean;
  signal type_cast_2927_inst_ack_1 : boolean;
  signal phi_stmt_2924_req_0 : boolean;
  signal phi_stmt_2911_ack_0 : boolean;
  signal phi_stmt_2918_ack_0 : boolean;
  signal phi_stmt_2924_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6792_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6792_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6792_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6792_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6792: Block -- control-path 
    signal convTransposeD_CP_6792_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6792_elements(0) <= convTransposeD_CP_6792_start;
    convTransposeD_CP_6792_symbol <= convTransposeD_CP_6792_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2591/$entry
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652__entry__
      -- CP-element group 0: 	 branch_block_stmt_2591/branch_block_stmt_2591__entry__
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_sample_start_
      -- 
    rr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(0), ack => RPIPE_Block3_start_2593_inst_req_0); -- 
    cr_6985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(0), ack => type_cast_2624_inst_req_1); -- 
    cr_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(0), ack => type_cast_2637_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2591/assign_stmt_2936__exit__
      -- CP-element group 1: 	 branch_block_stmt_2591/assign_stmt_2936__entry__
      -- CP-element group 1: 	 branch_block_stmt_2591/merge_stmt_2910__exit__
      -- CP-element group 1: 	 branch_block_stmt_2591/assign_stmt_2936/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/assign_stmt_2936/$exit
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Update/cr
      -- 
    rr_7513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2713_inst_req_0); -- 
    cr_7518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2713_inst_req_1); -- 
    rr_7536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2720_inst_req_0); -- 
    cr_7541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2720_inst_req_1); -- 
    rr_7559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2727_inst_req_0); -- 
    cr_7564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2727_inst_req_1); -- 
    rr_7582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2733_inst_req_0); -- 
    cr_7587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(1), ack => type_cast_2733_inst_req_1); -- 
    convTransposeD_CP_6792_elements(1) <= convTransposeD_CP_6792_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_update_start_
      -- 
    ra_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2593_inst_ack_0, ack => convTransposeD_CP_6792_elements(2)); -- 
    cr_6845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(2), ack => RPIPE_Block3_start_2593_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2593_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Sample/rr
      -- 
    ca_6846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2593_inst_ack_1, ack => convTransposeD_CP_6792_elements(3)); -- 
    rr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(3), ack => RPIPE_Block3_start_2596_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_update_start_
      -- 
    ra_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2596_inst_ack_0, ack => convTransposeD_CP_6792_elements(4)); -- 
    cr_6859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(4), ack => RPIPE_Block3_start_2596_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2596_Update/ca
      -- 
    ca_6860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2596_inst_ack_1, ack => convTransposeD_CP_6792_elements(5)); -- 
    rr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(5), ack => RPIPE_Block3_start_2599_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Sample/$exit
      -- 
    ra_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2599_inst_ack_0, ack => convTransposeD_CP_6792_elements(6)); -- 
    cr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(6), ack => RPIPE_Block3_start_2599_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2599_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Sample/rr
      -- 
    ca_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2599_inst_ack_1, ack => convTransposeD_CP_6792_elements(7)); -- 
    rr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(7), ack => RPIPE_Block3_start_2602_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Sample/ra
      -- 
    ra_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2602_inst_ack_0, ack => convTransposeD_CP_6792_elements(8)); -- 
    cr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(8), ack => RPIPE_Block3_start_2602_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2602_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_sample_start_
      -- 
    ca_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2602_inst_ack_1, ack => convTransposeD_CP_6792_elements(9)); -- 
    rr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(9), ack => RPIPE_Block3_start_2605_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Update/cr
      -- 
    ra_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2605_inst_ack_0, ack => convTransposeD_CP_6792_elements(10)); -- 
    cr_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(10), ack => RPIPE_Block3_start_2605_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2605_Update/$exit
      -- 
    ca_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2605_inst_ack_1, ack => convTransposeD_CP_6792_elements(11)); -- 
    rr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(11), ack => RPIPE_Block3_start_2608_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Sample/ra
      -- 
    ra_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2608_inst_ack_0, ack => convTransposeD_CP_6792_elements(12)); -- 
    cr_6915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(12), ack => RPIPE_Block3_start_2608_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2608_Update/$exit
      -- 
    ca_6916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2608_inst_ack_1, ack => convTransposeD_CP_6792_elements(13)); -- 
    rr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(13), ack => RPIPE_Block3_start_2611_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_sample_completed_
      -- 
    ra_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2611_inst_ack_0, ack => convTransposeD_CP_6792_elements(14)); -- 
    cr_6929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(14), ack => RPIPE_Block3_start_2611_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2611_update_completed_
      -- 
    ca_6930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2611_inst_ack_1, ack => convTransposeD_CP_6792_elements(15)); -- 
    rr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(15), ack => RPIPE_Block3_start_2614_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_update_start_
      -- 
    ra_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2614_inst_ack_0, ack => convTransposeD_CP_6792_elements(16)); -- 
    cr_6943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(16), ack => RPIPE_Block3_start_2614_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2614_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_sample_start_
      -- 
    ca_6944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2614_inst_ack_1, ack => convTransposeD_CP_6792_elements(17)); -- 
    rr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(17), ack => RPIPE_Block3_start_2617_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Sample/$exit
      -- 
    ra_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2617_inst_ack_0, ack => convTransposeD_CP_6792_elements(18)); -- 
    cr_6957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(18), ack => RPIPE_Block3_start_2617_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2617_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Sample/$entry
      -- 
    ca_6958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2617_inst_ack_1, ack => convTransposeD_CP_6792_elements(19)); -- 
    rr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(19), ack => RPIPE_Block3_start_2620_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_update_start_
      -- 
    ra_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2620_inst_ack_0, ack => convTransposeD_CP_6792_elements(20)); -- 
    cr_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(20), ack => RPIPE_Block3_start_2620_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2620_update_completed_
      -- 
    ca_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2620_inst_ack_1, ack => convTransposeD_CP_6792_elements(21)); -- 
    rr_6980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(21), ack => type_cast_2624_inst_req_0); -- 
    rr_6994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(21), ack => RPIPE_Block3_start_2633_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Sample/ra
      -- 
    ra_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2624_inst_ack_0, ack => convTransposeD_CP_6792_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2624_Update/ca
      -- 
    ca_6986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2624_inst_ack_1, ack => convTransposeD_CP_6792_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_update_start_
      -- 
    ra_6995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2633_inst_ack_0, ack => convTransposeD_CP_6792_elements(24)); -- 
    cr_6999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(24), ack => RPIPE_Block3_start_2633_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2633_update_completed_
      -- 
    ca_7000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2633_inst_ack_1, ack => convTransposeD_CP_6792_elements(25)); -- 
    rr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(25), ack => type_cast_2637_inst_req_0); -- 
    rr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(25), ack => RPIPE_Block3_start_2645_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Sample/$exit
      -- 
    ra_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2637_inst_ack_0, ack => convTransposeD_CP_6792_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/type_cast_2637_update_completed_
      -- 
    ca_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2637_inst_ack_1, ack => convTransposeD_CP_6792_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Update/cr
      -- 
    ra_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2645_inst_ack_0, ack => convTransposeD_CP_6792_elements(28)); -- 
    cr_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(28), ack => RPIPE_Block3_start_2645_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2645_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Sample/rr
      -- 
    ca_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2645_inst_ack_1, ack => convTransposeD_CP_6792_elements(29)); -- 
    rr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(29), ack => RPIPE_Block3_start_2648_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_update_start_
      -- 
    ra_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2648_inst_ack_0, ack => convTransposeD_CP_6792_elements(30)); -- 
    cr_7041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(30), ack => RPIPE_Block3_start_2648_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2648_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Sample/rr
      -- 
    ca_7042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2648_inst_ack_1, ack => convTransposeD_CP_6792_elements(31)); -- 
    rr_7050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(31), ack => RPIPE_Block3_start_2651_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Update/cr
      -- 
    ra_7051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2651_inst_ack_0, ack => convTransposeD_CP_6792_elements(32)); -- 
    cr_7055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(32), ack => RPIPE_Block3_start_2651_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/RPIPE_Block3_start_2651_Update/$exit
      -- 
    ca_7056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2651_inst_ack_1, ack => convTransposeD_CP_6792_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704__entry__
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/$entry
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652/$exit
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2594_to_assign_stmt_2652__exit__
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Update/$entry
      -- 
    cr_7072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2695_inst_req_1); -- 
    rr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2695_inst_req_0); -- 
    rr_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2699_inst_req_0); -- 
    rr_7095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2703_inst_req_0); -- 
    cr_7100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2703_inst_req_1); -- 
    cr_7086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(34), ack => type_cast_2699_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(23) & convTransposeD_CP_6792_elements(27) & convTransposeD_CP_6792_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Sample/$exit
      -- 
    ra_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_0, ack => convTransposeD_CP_6792_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2695_update_completed_
      -- 
    ca_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_1, ack => convTransposeD_CP_6792_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_sample_completed_
      -- 
    ra_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2699_inst_ack_0, ack => convTransposeD_CP_6792_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2699_Update/$exit
      -- 
    ca_7087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2699_inst_ack_1, ack => convTransposeD_CP_6792_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Sample/ra
      -- 
    ra_7096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2703_inst_ack_0, ack => convTransposeD_CP_6792_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/type_cast_2703_Update/ca
      -- 
    ca_7101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2703_inst_ack_1, ack => convTransposeD_CP_6792_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704__exit__
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2591/assign_stmt_2659_to_assign_stmt_2704/$exit
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2707/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2714/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2721/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Update/cr
      -- 
    rr_7487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(41), ack => type_cast_2731_inst_req_0); -- 
    cr_7492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(41), ack => type_cast_2731_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(36) & convTransposeD_CP_6792_elements(38) & convTransposeD_CP_6792_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Sample/$exit
      -- 
    ra_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2768_inst_ack_0, ack => convTransposeD_CP_6792_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Update/$exit
      -- 
    ca_7118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2768_inst_ack_1, ack => convTransposeD_CP_6792_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Sample/ra
      -- 
    ra_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_0, ack => convTransposeD_CP_6792_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Update/$exit
      -- 
    ca_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_1, ack => convTransposeD_CP_6792_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Sample/ra
      -- 
    ra_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2776_inst_ack_0, ack => convTransposeD_CP_6792_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Update/$exit
      -- 
    ca_7146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2776_inst_ack_1, ack => convTransposeD_CP_6792_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Sample/ra
      -- 
    ra_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2806_inst_ack_0, ack => convTransposeD_CP_6792_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_index_scale_1/scale_rename_ack
      -- 
    ca_7160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2806_inst_ack_1, ack => convTransposeD_CP_6792_elements(49)); -- 
    req_7185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(49), ack => array_obj_ref_2812_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_sample_complete
      -- 
    ack_7186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2812_index_offset_ack_0, ack => convTransposeD_CP_6792_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_request/req
      -- 
    ack_7191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2812_index_offset_ack_1, ack => convTransposeD_CP_6792_elements(51)); -- 
    req_7200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(51), ack => addr_of_2813_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_request/ack
      -- 
    ack_7201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2813_final_reg_ack_0, ack => convTransposeD_CP_6792_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/word_access_start/word_0/rr
      -- 
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2813_final_reg_ack_1, ack => convTransposeD_CP_6792_elements(53)); -- 
    rr_7239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(53), ack => ptr_deref_2817_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Sample/word_access_start/word_0/ra
      -- 
    ra_7240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2817_load_0_ack_0, ack => convTransposeD_CP_6792_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/ptr_deref_2817_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/ptr_deref_2817_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/ptr_deref_2817_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/ptr_deref_2817_Merge/merge_ack
      -- 
    ca_7251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2817_load_0_ack_1, ack => convTransposeD_CP_6792_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Sample/req
      -- 
    req_7281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(56), ack => array_obj_ref_2835_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(43) & convTransposeD_CP_6792_elements(45) & convTransposeD_CP_6792_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Sample/ack
      -- 
    ack_7282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2835_index_offset_ack_0, ack => convTransposeD_CP_6792_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_request/req
      -- 
    ack_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2835_index_offset_ack_1, ack => convTransposeD_CP_6792_elements(58)); -- 
    req_7296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(58), ack => addr_of_2836_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_request/ack
      -- 
    ack_7297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2836_final_reg_ack_0, ack => convTransposeD_CP_6792_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_word_addrgen/root_register_ack
      -- 
    ack_7302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2836_final_reg_ack_1, ack => convTransposeD_CP_6792_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/ptr_deref_2839_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/ptr_deref_2839_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/ptr_deref_2839_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/ptr_deref_2839_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/word_access_start/word_0/rr
      -- 
    rr_7340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(61), ack => ptr_deref_2839_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(55) & convTransposeD_CP_6792_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Sample/word_access_start/word_0/ra
      -- 
    ra_7341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2839_store_0_ack_0, ack => convTransposeD_CP_6792_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/word_access_complete/word_0/ca
      -- 
    ca_7352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2839_store_0_ack_1, ack => convTransposeD_CP_6792_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Sample/ra
      -- 
    ra_7361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2844_inst_ack_0, ack => convTransposeD_CP_6792_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Update/ca
      -- 
    ca_7366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2844_inst_ack_1, ack => convTransposeD_CP_6792_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857__entry__
      -- CP-element group 66: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856__exit__
      -- CP-element group 66: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/$exit
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2591/R_cmp_2858_place
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2591/if_stmt_2857_else_link/$entry
      -- 
    branch_req_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(66), ack => if_stmt_2857_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(50) & convTransposeD_CP_6792_elements(57) & convTransposeD_CP_6792_elements(63) & convTransposeD_CP_6792_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2591/merge_stmt_2863__exit__
      -- CP-element group 67: 	 branch_block_stmt_2591/assign_stmt_2869__entry__
      -- CP-element group 67: 	 branch_block_stmt_2591/assign_stmt_2869__exit__
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2591/if_stmt_2857_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2591/if_stmt_2857_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2591/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2591/assign_stmt_2869/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/assign_stmt_2869/$exit
      -- CP-element group 67: 	 branch_block_stmt_2591/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2591/merge_stmt_2863_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2591/merge_stmt_2863_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/merge_stmt_2863_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2591/merge_stmt_2863_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2857_branch_ack_1, ack => convTransposeD_CP_6792_elements(67)); -- 
    rr_7697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2914_inst_req_0); -- 
    cr_7702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2914_inst_req_1); -- 
    rr_7720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2921_inst_req_0); -- 
    cr_7725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2921_inst_req_1); -- 
    rr_7743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2927_inst_req_0); -- 
    cr_7748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(67), ack => type_cast_2927_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2591/merge_stmt_2871__exit__
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903__entry__
      -- CP-element group 68: 	 branch_block_stmt_2591/if_stmt_2857_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2591/if_stmt_2857_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2591/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/$entry
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2591/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2591/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2591/merge_stmt_2871_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2591/merge_stmt_2871_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2591/merge_stmt_2871_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2591/merge_stmt_2871_PhiAck/dummy
      -- 
    else_choice_transition_7383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2857_branch_ack_0, ack => convTransposeD_CP_6792_elements(68)); -- 
    rr_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(68), ack => type_cast_2885_inst_req_0); -- 
    cr_7404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(68), ack => type_cast_2885_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Sample/ra
      -- 
    ra_7400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2885_inst_ack_0, ack => convTransposeD_CP_6792_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904__entry__
      -- CP-element group 70: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903__exit__
      -- CP-element group 70: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/$exit
      -- CP-element group 70: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2591/assign_stmt_2877_to_assign_stmt_2903/type_cast_2885_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2591/R_cmp121_2905_place
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2591/if_stmt_2904_else_link/$entry
      -- 
    ca_7405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2885_inst_ack_1, ack => convTransposeD_CP_6792_elements(70)); -- 
    branch_req_7413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(70), ack => if_stmt_2904_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2591/assign_stmt_2943__entry__
      -- CP-element group 71: 	 branch_block_stmt_2591/merge_stmt_2938__exit__
      -- CP-element group 71: 	 branch_block_stmt_2591/if_stmt_2904_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2591/if_stmt_2904_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2591/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2591/assign_stmt_2943/$entry
      -- CP-element group 71: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2591/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2591/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2591/merge_stmt_2938_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2591/merge_stmt_2938_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2591/merge_stmt_2938_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2591/merge_stmt_2938_PhiAck/dummy
      -- 
    if_choice_transition_7418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2904_branch_ack_1, ack => convTransposeD_CP_6792_elements(71)); -- 
    req_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(71), ack => WPIPE_Block3_done_2940_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2591/if_stmt_2904_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2591/if_stmt_2904_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2911/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2904_branch_ack_0, ack => convTransposeD_CP_6792_elements(72)); -- 
    rr_7648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2923_inst_req_0); -- 
    cr_7653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2923_inst_req_1); -- 
    rr_7671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2929_inst_req_0); -- 
    cr_7676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(72), ack => type_cast_2929_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Update/req
      -- 
    ack_7439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2940_inst_ack_0, ack => convTransposeD_CP_6792_elements(73)); -- 
    req_7443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(73), ack => WPIPE_Block3_done_2940_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2591/branch_block_stmt_2591__exit__
      -- CP-element group 74: 	 branch_block_stmt_2591/assign_stmt_2943__exit__
      -- CP-element group 74: 	 branch_block_stmt_2591/$exit
      -- CP-element group 74: 	 branch_block_stmt_2591/return__
      -- CP-element group 74: 	 branch_block_stmt_2591/merge_stmt_2945__exit__
      -- CP-element group 74: 	 branch_block_stmt_2591/assign_stmt_2943/$exit
      -- CP-element group 74: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2591/assign_stmt_2943/WPIPE_Block3_done_2940_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2591/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2591/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2591/merge_stmt_2945_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2591/merge_stmt_2945_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2591/merge_stmt_2945_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2591/merge_stmt_2945_PhiAck/dummy
      -- 
    ack_7444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2940_inst_ack_1, ack => convTransposeD_CP_6792_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2707/$exit
      -- CP-element group 75: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2711_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_req
      -- 
    phi_stmt_2707_req_7455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2707_req_7455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(75), ack => phi_stmt_2707_req_0); -- 
    -- Element group convTransposeD_CP_6792_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(41), ack => convTransposeD_CP_6792_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2714/$exit
      -- CP-element group 76: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2718_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_req
      -- 
    phi_stmt_2714_req_7463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2714_req_7463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(76), ack => phi_stmt_2714_req_0); -- 
    -- Element group convTransposeD_CP_6792_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(41), ack => convTransposeD_CP_6792_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2721/$exit
      -- CP-element group 77: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2725_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_req
      -- 
    phi_stmt_2721_req_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2721_req_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(77), ack => phi_stmt_2721_req_0); -- 
    -- Element group convTransposeD_CP_6792_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(41), ack => convTransposeD_CP_6792_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Sample/ra
      -- 
    ra_7488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2731_inst_ack_0, ack => convTransposeD_CP_6792_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/Update/ca
      -- 
    ca_7493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2731_inst_ack_1, ack => convTransposeD_CP_6792_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/$exit
      -- CP-element group 80: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/$exit
      -- CP-element group 80: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2731/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_req
      -- 
    phi_stmt_2728_req_7494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2728_req_7494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(80), ack => phi_stmt_2728_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(78) & convTransposeD_CP_6792_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2591/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(75) & convTransposeD_CP_6792_elements(76) & convTransposeD_CP_6792_elements(77) & convTransposeD_CP_6792_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Sample/ra
      -- 
    ra_7514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_0, ack => convTransposeD_CP_6792_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/Update/ca
      -- 
    ca_7519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_1, ack => convTransposeD_CP_6792_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/$exit
      -- CP-element group 84: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/$exit
      -- CP-element group 84: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_sources/type_cast_2713/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2707/phi_stmt_2707_req
      -- 
    phi_stmt_2707_req_7520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2707_req_7520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(84), ack => phi_stmt_2707_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(82) & convTransposeD_CP_6792_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Sample/ra
      -- 
    ra_7537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2720_inst_ack_0, ack => convTransposeD_CP_6792_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/Update/ca
      -- 
    ca_7542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2720_inst_ack_1, ack => convTransposeD_CP_6792_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/$exit
      -- CP-element group 87: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/$exit
      -- CP-element group 87: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_sources/type_cast_2720/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2714/phi_stmt_2714_req
      -- 
    phi_stmt_2714_req_7543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2714_req_7543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(87), ack => phi_stmt_2714_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(85) & convTransposeD_CP_6792_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Sample/ra
      -- 
    ra_7560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2727_inst_ack_0, ack => convTransposeD_CP_6792_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/Update/ca
      -- 
    ca_7565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2727_inst_ack_1, ack => convTransposeD_CP_6792_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/$exit
      -- CP-element group 90: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/$exit
      -- CP-element group 90: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_sources/type_cast_2727/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2721/phi_stmt_2721_req
      -- 
    phi_stmt_2721_req_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2721_req_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(90), ack => phi_stmt_2721_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(88) & convTransposeD_CP_6792_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Sample/ra
      -- 
    ra_7583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2733_inst_ack_0, ack => convTransposeD_CP_6792_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/Update/ca
      -- 
    ca_7588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2733_inst_ack_1, ack => convTransposeD_CP_6792_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/$exit
      -- CP-element group 93: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/$exit
      -- CP-element group 93: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_sources/type_cast_2733/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2728/phi_stmt_2728_req
      -- 
    phi_stmt_2728_req_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2728_req_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(93), ack => phi_stmt_2728_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(91) & convTransposeD_CP_6792_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2591/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(84) & convTransposeD_CP_6792_elements(87) & convTransposeD_CP_6792_elements(90) & convTransposeD_CP_6792_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2591/merge_stmt_2706_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2591/merge_stmt_2706_PhiAck/$entry
      -- 
    convTransposeD_CP_6792_elements(95) <= OrReduce(convTransposeD_CP_6792_elements(81) & convTransposeD_CP_6792_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2591/merge_stmt_2706_PhiAck/phi_stmt_2707_ack
      -- 
    phi_stmt_2707_ack_7594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2707_ack_0, ack => convTransposeD_CP_6792_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2591/merge_stmt_2706_PhiAck/phi_stmt_2714_ack
      -- 
    phi_stmt_2714_ack_7595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2714_ack_0, ack => convTransposeD_CP_6792_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2591/merge_stmt_2706_PhiAck/phi_stmt_2721_ack
      -- 
    phi_stmt_2721_ack_7596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2721_ack_0, ack => convTransposeD_CP_6792_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2591/merge_stmt_2706_PhiAck/phi_stmt_2728_ack
      -- 
    phi_stmt_2728_ack_7597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2728_ack_0, ack => convTransposeD_CP_6792_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856__entry__
      -- CP-element group 100: 	 branch_block_stmt_2591/merge_stmt_2706__exit__
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2812_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2813_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2806_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2768_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2776_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2772_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2817_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/array_obj_ref_2835_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/addr_of_2836_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/ptr_deref_2839_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2591/assign_stmt_2740_to_assign_stmt_2856/type_cast_2844_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2591/merge_stmt_2706_PhiAck/$exit
      -- 
    rr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2768_inst_req_0); -- 
    cr_7159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2806_inst_req_1); -- 
    cr_7117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2768_inst_req_1); -- 
    req_7190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => array_obj_ref_2812_index_offset_req_1); -- 
    cr_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2776_inst_req_1); -- 
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => addr_of_2813_final_reg_req_1); -- 
    rr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2806_inst_req_0); -- 
    rr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2772_inst_req_0); -- 
    rr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2776_inst_req_0); -- 
    cr_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2772_inst_req_1); -- 
    cr_7250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => ptr_deref_2817_load_0_req_1); -- 
    req_7286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => array_obj_ref_2835_index_offset_req_1); -- 
    req_7301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => addr_of_2836_final_reg_req_1); -- 
    cr_7351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => ptr_deref_2839_store_0_req_1); -- 
    rr_7360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2844_inst_req_0); -- 
    cr_7365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(100), ack => type_cast_2844_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(96) & convTransposeD_CP_6792_elements(97) & convTransposeD_CP_6792_elements(98) & convTransposeD_CP_6792_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2911/$exit
      -- CP-element group 101: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2917_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_req
      -- 
    phi_stmt_2911_req_7632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2911_req_7632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(101), ack => phi_stmt_2911_req_1); -- 
    -- Element group convTransposeD_CP_6792_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6792_elements(72), ack => convTransposeD_CP_6792_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Sample/ra
      -- 
    ra_7649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_0, ack => convTransposeD_CP_6792_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/Update/ca
      -- 
    ca_7654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_1, ack => convTransposeD_CP_6792_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/$exit
      -- CP-element group 104: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/$exit
      -- CP-element group 104: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2923/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_req
      -- 
    phi_stmt_2918_req_7655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2918_req_7655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(104), ack => phi_stmt_2918_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(102) & convTransposeD_CP_6792_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Sample/ra
      -- 
    ra_7672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2929_inst_ack_0, ack => convTransposeD_CP_6792_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/Update/ca
      -- 
    ca_7677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2929_inst_ack_1, ack => convTransposeD_CP_6792_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/$exit
      -- CP-element group 107: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/$exit
      -- CP-element group 107: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2929/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_req
      -- 
    phi_stmt_2924_req_7678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2924_req_7678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(107), ack => phi_stmt_2924_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(105) & convTransposeD_CP_6792_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2591/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(101) & convTransposeD_CP_6792_elements(104) & convTransposeD_CP_6792_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Sample/ra
      -- 
    ra_7698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_0, ack => convTransposeD_CP_6792_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/Update/ca
      -- 
    ca_7703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_1, ack => convTransposeD_CP_6792_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/$exit
      -- CP-element group 111: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/$exit
      -- CP-element group 111: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_sources/type_cast_2914/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2911/phi_stmt_2911_req
      -- 
    phi_stmt_2911_req_7704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2911_req_7704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(111), ack => phi_stmt_2911_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(109) & convTransposeD_CP_6792_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Sample/ra
      -- 
    ra_7721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2921_inst_ack_0, ack => convTransposeD_CP_6792_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/Update/ca
      -- 
    ca_7726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2921_inst_ack_1, ack => convTransposeD_CP_6792_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/$exit
      -- CP-element group 114: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/$exit
      -- CP-element group 114: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_sources/type_cast_2921/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2918/phi_stmt_2918_req
      -- 
    phi_stmt_2918_req_7727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2918_req_7727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(114), ack => phi_stmt_2918_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(112) & convTransposeD_CP_6792_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Sample/ra
      -- 
    ra_7744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2927_inst_ack_0, ack => convTransposeD_CP_6792_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/Update/ca
      -- 
    ca_7749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2927_inst_ack_1, ack => convTransposeD_CP_6792_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/$exit
      -- CP-element group 117: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/$exit
      -- CP-element group 117: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_sources/type_cast_2927/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2924/phi_stmt_2924_req
      -- 
    phi_stmt_2924_req_7750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2924_req_7750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6792_elements(117), ack => phi_stmt_2924_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(115) & convTransposeD_CP_6792_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2591/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(111) & convTransposeD_CP_6792_elements(114) & convTransposeD_CP_6792_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2591/merge_stmt_2910_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2591/merge_stmt_2910_PhiAck/$entry
      -- 
    convTransposeD_CP_6792_elements(119) <= OrReduce(convTransposeD_CP_6792_elements(108) & convTransposeD_CP_6792_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2591/merge_stmt_2910_PhiAck/phi_stmt_2911_ack
      -- 
    phi_stmt_2911_ack_7755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2911_ack_0, ack => convTransposeD_CP_6792_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2591/merge_stmt_2910_PhiAck/phi_stmt_2918_ack
      -- 
    phi_stmt_2918_ack_7756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2918_ack_0, ack => convTransposeD_CP_6792_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2591/merge_stmt_2910_PhiAck/phi_stmt_2924_ack
      -- 
    phi_stmt_2924_ack_7757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2924_ack_0, ack => convTransposeD_CP_6792_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2591/merge_stmt_2910_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6792_elements(120) & convTransposeD_CP_6792_elements(121) & convTransposeD_CP_6792_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6792_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2834_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2834_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2811_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2811_scaled : std_logic_vector(13 downto 0);
    signal add103_2869 : std_logic_vector(15 downto 0);
    signal add32_2670 : std_logic_vector(15 downto 0);
    signal add50_2676 : std_logic_vector(15 downto 0);
    signal add63_2687 : std_logic_vector(15 downto 0);
    signal add82_2787 : std_logic_vector(63 downto 0);
    signal add84_2797 : std_logic_vector(63 downto 0);
    signal add96_2851 : std_logic_vector(31 downto 0);
    signal add_2643 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2745 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2812_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2812_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2812_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2812_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2812_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2812_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2835_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2835_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2835_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2835_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2835_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2835_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2814 : std_logic_vector(31 downto 0);
    signal arrayidx92_2837 : std_logic_vector(31 downto 0);
    signal call11_2612 : std_logic_vector(15 downto 0);
    signal call13_2615 : std_logic_vector(15 downto 0);
    signal call14_2618 : std_logic_vector(15 downto 0);
    signal call15_2621 : std_logic_vector(15 downto 0);
    signal call16_2634 : std_logic_vector(15 downto 0);
    signal call18_2646 : std_logic_vector(15 downto 0);
    signal call1_2597 : std_logic_vector(15 downto 0);
    signal call20_2649 : std_logic_vector(15 downto 0);
    signal call22_2652 : std_logic_vector(15 downto 0);
    signal call3_2600 : std_logic_vector(15 downto 0);
    signal call5_2603 : std_logic_vector(15 downto 0);
    signal call7_2606 : std_logic_vector(15 downto 0);
    signal call9_2609 : std_logic_vector(15 downto 0);
    signal call_2594 : std_logic_vector(15 downto 0);
    signal cmp111_2882 : std_logic_vector(0 downto 0);
    signal cmp121_2903 : std_logic_vector(0 downto 0);
    signal cmp_2856 : std_logic_vector(0 downto 0);
    signal conv17_2638 : std_logic_vector(31 downto 0);
    signal conv70_2769 : std_logic_vector(63 downto 0);
    signal conv73_2696 : std_logic_vector(63 downto 0);
    signal conv75_2773 : std_logic_vector(63 downto 0);
    signal conv78_2700 : std_logic_vector(63 downto 0);
    signal conv80_2777 : std_logic_vector(63 downto 0);
    signal conv95_2845 : std_logic_vector(31 downto 0);
    signal conv99_2704 : std_logic_vector(31 downto 0);
    signal conv_2625 : std_logic_vector(31 downto 0);
    signal idxprom91_2830 : std_logic_vector(63 downto 0);
    signal idxprom_2807 : std_logic_vector(63 downto 0);
    signal inc115_2886 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2891 : std_logic_vector(15 downto 0);
    signal inc_2877 : std_logic_vector(15 downto 0);
    signal indvar_2707 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2936 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2924 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2728 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2918 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2721 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2898 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2911 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2714 : std_logic_vector(15 downto 0);
    signal mul59_2760 : std_logic_vector(15 downto 0);
    signal mul81_2782 : std_logic_vector(63 downto 0);
    signal mul83_2792 : std_logic_vector(63 downto 0);
    signal mul_2750 : std_logic_vector(15 downto 0);
    signal ptr_deref_2817_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2817_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2817_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2817_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2817_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2839_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2839_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2839_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2839_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2839_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2839_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2631 : std_logic_vector(31 downto 0);
    signal shr135_2659 : std_logic_vector(15 downto 0);
    signal shr31136_2665 : std_logic_vector(15 downto 0);
    signal shr86_2803 : std_logic_vector(31 downto 0);
    signal shr90_2824 : std_logic_vector(63 downto 0);
    signal sub53_2755 : std_logic_vector(15 downto 0);
    signal sub66_2692 : std_logic_vector(15 downto 0);
    signal sub67_2765 : std_logic_vector(15 downto 0);
    signal sub_2681 : std_logic_vector(15 downto 0);
    signal tmp1_2740 : std_logic_vector(31 downto 0);
    signal tmp88_2818 : std_logic_vector(63 downto 0);
    signal type_cast_2629_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2657_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2663_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2674_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2685_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2711_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2713_wire : std_logic_vector(31 downto 0);
    signal type_cast_2718_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2720_wire : std_logic_vector(15 downto 0);
    signal type_cast_2725_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2727_wire : std_logic_vector(15 downto 0);
    signal type_cast_2731_wire : std_logic_vector(15 downto 0);
    signal type_cast_2733_wire : std_logic_vector(15 downto 0);
    signal type_cast_2738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2801_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2822_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2828_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2849_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2867_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2875_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2895_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2914_wire : std_logic_vector(15 downto 0);
    signal type_cast_2917_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2921_wire : std_logic_vector(15 downto 0);
    signal type_cast_2923_wire : std_logic_vector(15 downto 0);
    signal type_cast_2927_wire : std_logic_vector(15 downto 0);
    signal type_cast_2929_wire : std_logic_vector(15 downto 0);
    signal type_cast_2934_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2942_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2812_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2812_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2812_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2812_resized_base_address <= "00000000000000";
    array_obj_ref_2835_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2835_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2835_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2835_resized_base_address <= "00000000000000";
    ptr_deref_2817_word_offset_0 <= "00000000000000";
    ptr_deref_2839_word_offset_0 <= "00000000000000";
    type_cast_2629_wire_constant <= "00000000000000000000000000010000";
    type_cast_2657_wire_constant <= "0000000000000010";
    type_cast_2663_wire_constant <= "0000000000000001";
    type_cast_2674_wire_constant <= "1111111111111111";
    type_cast_2685_wire_constant <= "1111111111111111";
    type_cast_2711_wire_constant <= "00000000000000000000000000000000";
    type_cast_2718_wire_constant <= "0000000000000000";
    type_cast_2725_wire_constant <= "0000000000000000";
    type_cast_2738_wire_constant <= "00000000000000000000000000000100";
    type_cast_2801_wire_constant <= "00000000000000000000000000000010";
    type_cast_2822_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2828_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2849_wire_constant <= "00000000000000000000000000000100";
    type_cast_2867_wire_constant <= "0000000000000100";
    type_cast_2875_wire_constant <= "0000000000000001";
    type_cast_2895_wire_constant <= "0000000000000000";
    type_cast_2917_wire_constant <= "0000000000000000";
    type_cast_2934_wire_constant <= "00000000000000000000000000000001";
    type_cast_2942_wire_constant <= "0000000000000001";
    phi_stmt_2707: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2711_wire_constant & type_cast_2713_wire;
      req <= phi_stmt_2707_req_0 & phi_stmt_2707_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2707",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2707_ack_0,
          idata => idata,
          odata => indvar_2707,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2707
    phi_stmt_2714: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2718_wire_constant & type_cast_2720_wire;
      req <= phi_stmt_2714_req_0 & phi_stmt_2714_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2714",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2714_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2714,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2714
    phi_stmt_2721: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2725_wire_constant & type_cast_2727_wire;
      req <= phi_stmt_2721_req_0 & phi_stmt_2721_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2721",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2721_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2721,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2721
    phi_stmt_2728: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2731_wire & type_cast_2733_wire;
      req <= phi_stmt_2728_req_0 & phi_stmt_2728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2728",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2728_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2728
    phi_stmt_2911: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2914_wire & type_cast_2917_wire_constant;
      req <= phi_stmt_2911_req_0 & phi_stmt_2911_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2911",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2911_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2911,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2911
    phi_stmt_2918: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2921_wire & type_cast_2923_wire;
      req <= phi_stmt_2918_req_0 & phi_stmt_2918_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2918",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2918_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2918,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2918
    phi_stmt_2924: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2927_wire & type_cast_2929_wire;
      req <= phi_stmt_2924_req_0 & phi_stmt_2924_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2924",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2924_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2924,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2924
    -- flow-through select operator MUX_2897_inst
    input_dim1x_x2_2898 <= type_cast_2895_wire_constant when (cmp111_2882(0) /=  '0') else inc_2877;
    addr_of_2813_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2813_final_reg_req_0;
      addr_of_2813_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2813_final_reg_req_1;
      addr_of_2813_final_reg_ack_1<= rack(0);
      addr_of_2813_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2813_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2812_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2836_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2836_final_reg_req_0;
      addr_of_2836_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2836_final_reg_req_1;
      addr_of_2836_final_reg_ack_1<= rack(0);
      addr_of_2836_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2836_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2835_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2837,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2624_inst_req_0;
      type_cast_2624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2624_inst_req_1;
      type_cast_2624_inst_ack_1<= rack(0);
      type_cast_2624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2637_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2637_inst_req_0;
      type_cast_2637_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2637_inst_req_1;
      type_cast_2637_inst_ack_1<= rack(0);
      type_cast_2637_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2637_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2634,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2638,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2695_inst_req_0;
      type_cast_2695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2695_inst_req_1;
      type_cast_2695_inst_ack_1<= rack(0);
      type_cast_2695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2652,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2699_inst_req_0;
      type_cast_2699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2699_inst_req_1;
      type_cast_2699_inst_ack_1<= rack(0);
      type_cast_2699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2703_inst_req_0;
      type_cast_2703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2703_inst_req_1;
      type_cast_2703_inst_ack_1<= rack(0);
      type_cast_2703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2600,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2704,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2713_inst_req_0;
      type_cast_2713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2713_inst_req_1;
      type_cast_2713_inst_ack_1<= rack(0);
      type_cast_2713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2936,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2713_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2720_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2720_inst_req_0;
      type_cast_2720_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2720_inst_req_1;
      type_cast_2720_inst_ack_1<= rack(0);
      type_cast_2720_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2720_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2720_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2727_inst_req_0;
      type_cast_2727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2727_inst_req_1;
      type_cast_2727_inst_ack_1<= rack(0);
      type_cast_2727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2918,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2727_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2731_inst_req_0;
      type_cast_2731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2731_inst_req_1;
      type_cast_2731_inst_ack_1<= rack(0);
      type_cast_2731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2731_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2733_inst_req_0;
      type_cast_2733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2733_inst_req_1;
      type_cast_2733_inst_ack_1<= rack(0);
      type_cast_2733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2733_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2768_inst_req_0;
      type_cast_2768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2768_inst_req_1;
      type_cast_2768_inst_ack_1<= rack(0);
      type_cast_2768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2772_inst_req_0;
      type_cast_2772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2772_inst_req_1;
      type_cast_2772_inst_ack_1<= rack(0);
      type_cast_2772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2776_inst_req_0;
      type_cast_2776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2776_inst_req_1;
      type_cast_2776_inst_ack_1<= rack(0);
      type_cast_2776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2806_inst_req_0;
      type_cast_2806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2806_inst_req_1;
      type_cast_2806_inst_ack_1<= rack(0);
      type_cast_2806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2844_inst_req_0;
      type_cast_2844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2844_inst_req_1;
      type_cast_2844_inst_ack_1<= rack(0);
      type_cast_2844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2885_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2885_inst_req_0;
      type_cast_2885_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2885_inst_req_1;
      type_cast_2885_inst_ack_1<= rack(0);
      type_cast_2885_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2885_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2886,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2914_inst_req_0;
      type_cast_2914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2914_inst_req_1;
      type_cast_2914_inst_ack_1<= rack(0);
      type_cast_2914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2869,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2914_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2921_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2921_inst_req_0;
      type_cast_2921_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2921_inst_req_1;
      type_cast_2921_inst_ack_1<= rack(0);
      type_cast_2921_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2921_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2921_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2923_inst_req_0;
      type_cast_2923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2923_inst_req_1;
      type_cast_2923_inst_ack_1<= rack(0);
      type_cast_2923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2927_inst_req_0;
      type_cast_2927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2927_inst_req_1;
      type_cast_2927_inst_ack_1<= rack(0);
      type_cast_2927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2927_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2929_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2929_inst_req_0;
      type_cast_2929_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2929_inst_req_1;
      type_cast_2929_inst_ack_1<= rack(0);
      type_cast_2929_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2929_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2929_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2812_index_1_rename
    process(R_idxprom_2811_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2811_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2811_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2812_index_1_resize
    process(idxprom_2807) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2807;
      ov := iv(13 downto 0);
      R_idxprom_2811_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2812_root_address_inst
    process(array_obj_ref_2812_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2812_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2812_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2835_index_1_rename
    process(R_idxprom91_2834_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2834_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2834_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2835_index_1_resize
    process(idxprom91_2830) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2830;
      ov := iv(13 downto 0);
      R_idxprom91_2834_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2835_root_address_inst
    process(array_obj_ref_2835_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2835_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2835_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_addr_0
    process(ptr_deref_2817_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2817_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2817_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_base_resize
    process(arrayidx87_2814) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2814;
      ov := iv(13 downto 0);
      ptr_deref_2817_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_gather_scatter
    process(ptr_deref_2817_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2817_data_0;
      ov(63 downto 0) := iv;
      tmp88_2818 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_root_address_inst
    process(ptr_deref_2817_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2817_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2817_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2839_addr_0
    process(ptr_deref_2839_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2839_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2839_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2839_base_resize
    process(arrayidx92_2837) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2837;
      ov := iv(13 downto 0);
      ptr_deref_2839_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2839_gather_scatter
    process(tmp88_2818) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2818;
      ov(63 downto 0) := iv;
      ptr_deref_2839_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2839_root_address_inst
    process(ptr_deref_2839_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2839_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2839_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2857_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2856;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2857_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2857_branch_req_0,
          ack0 => if_stmt_2857_branch_ack_0,
          ack1 => if_stmt_2857_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2904_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2903;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2904_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2904_branch_req_0,
          ack0 => if_stmt_2904_branch_ack_0,
          ack1 => if_stmt_2904_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2669_inst
    process(shr135_2659, shr31136_2665) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2659, shr31136_2665, tmp_var);
      add32_2670 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2675_inst
    process(call7_2606) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2606, type_cast_2674_wire_constant, tmp_var);
      add50_2676 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2686_inst
    process(call9_2609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2609, type_cast_2685_wire_constant, tmp_var);
      add63_2687 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2754_inst
    process(sub_2681, mul_2750) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2681, mul_2750, tmp_var);
      sub53_2755 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2764_inst
    process(sub66_2692, mul59_2760) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2692, mul59_2760, tmp_var);
      sub67_2765 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2868_inst
    process(input_dim2x_x1_2714) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2714, type_cast_2867_wire_constant, tmp_var);
      add103_2869 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2876_inst
    process(input_dim1x_x1_2721) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2721, type_cast_2875_wire_constant, tmp_var);
      inc_2877 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2890_inst
    process(inc115_2886, input_dim0x_x2_2728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2886, input_dim0x_x2_2728, tmp_var);
      inc115x_xinput_dim0x_x2_2891 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2744_inst
    process(add_2643, tmp1_2740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2643, tmp1_2740, tmp_var);
      add_src_0x_x0_2745 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2850_inst
    process(conv95_2845) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2845, type_cast_2849_wire_constant, tmp_var);
      add96_2851 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2935_inst
    process(indvar_2707) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2707, type_cast_2934_wire_constant, tmp_var);
      indvarx_xnext_2936 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2786_inst
    process(mul81_2782, conv75_2773) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2782, conv75_2773, tmp_var);
      add82_2787 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2796_inst
    process(mul83_2792, conv70_2769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2792, conv70_2769, tmp_var);
      add84_2797 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2829_inst
    process(shr90_2824) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2824, type_cast_2828_wire_constant, tmp_var);
      idxprom91_2830 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2881_inst
    process(inc_2877, call1_2597) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2877, call1_2597, tmp_var);
      cmp111_2882 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2902_inst
    process(inc115x_xinput_dim0x_x2_2891, call_2594) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2891, call_2594, tmp_var);
      cmp121_2903 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2658_inst
    process(call_2594) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2594, type_cast_2657_wire_constant, tmp_var);
      shr135_2659 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2664_inst
    process(call_2594) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2594, type_cast_2663_wire_constant, tmp_var);
      shr31136_2665 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2802_inst
    process(add_src_0x_x0_2745) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2745, type_cast_2801_wire_constant, tmp_var);
      shr86_2803 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2823_inst
    process(add84_2797) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2797, type_cast_2822_wire_constant, tmp_var);
      shr90_2824 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2749_inst
    process(input_dim0x_x2_2728, call13_2615) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2728, call13_2615, tmp_var);
      mul_2750 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2759_inst
    process(input_dim1x_x1_2721, call13_2615) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2721, call13_2615, tmp_var);
      mul59_2760 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2739_inst
    process(indvar_2707) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2707, type_cast_2738_wire_constant, tmp_var);
      tmp1_2740 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2781_inst
    process(conv80_2777, conv78_2700) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2777, conv78_2700, tmp_var);
      mul81_2782 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2791_inst
    process(add82_2787, conv73_2696) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2787, conv73_2696, tmp_var);
      mul83_2792 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2642_inst
    process(shl_2631, conv17_2638) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2631, conv17_2638, tmp_var);
      add_2643 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2630_inst
    process(conv_2625) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2625, type_cast_2629_wire_constant, tmp_var);
      shl_2631 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2680_inst
    process(add50_2676, call14_2618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2676, call14_2618, tmp_var);
      sub_2681 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2691_inst
    process(add63_2687, call14_2618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2687, call14_2618, tmp_var);
      sub66_2692 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2855_inst
    process(add96_2851, conv99_2704) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2851, conv99_2704, tmp_var);
      cmp_2856 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2812_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2811_scaled;
      array_obj_ref_2812_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2812_index_offset_req_0;
      array_obj_ref_2812_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2812_index_offset_req_1;
      array_obj_ref_2812_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2835_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2834_scaled;
      array_obj_ref_2835_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2835_index_offset_req_0;
      array_obj_ref_2835_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2835_index_offset_req_1;
      array_obj_ref_2835_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2817_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2817_load_0_req_0;
      ptr_deref_2817_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2817_load_0_req_1;
      ptr_deref_2817_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2817_word_address_0;
      ptr_deref_2817_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2839_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2839_store_0_req_0;
      ptr_deref_2839_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2839_store_0_req_1;
      ptr_deref_2839_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2839_word_address_0;
      data_in <= ptr_deref_2839_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2593_inst RPIPE_Block3_start_2596_inst RPIPE_Block3_start_2599_inst RPIPE_Block3_start_2602_inst RPIPE_Block3_start_2605_inst RPIPE_Block3_start_2608_inst RPIPE_Block3_start_2611_inst RPIPE_Block3_start_2614_inst RPIPE_Block3_start_2617_inst RPIPE_Block3_start_2620_inst RPIPE_Block3_start_2633_inst RPIPE_Block3_start_2645_inst RPIPE_Block3_start_2648_inst RPIPE_Block3_start_2651_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2593_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2596_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2599_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2602_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2605_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2608_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2611_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2614_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2617_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2620_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2633_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2645_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2648_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2651_inst_req_0;
      RPIPE_Block3_start_2593_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2596_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2599_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2602_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2605_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2608_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2611_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2614_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2617_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2620_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2633_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2645_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2648_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2651_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2593_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2596_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2599_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2602_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2605_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2608_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2611_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2614_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2617_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2620_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2633_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2645_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2648_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2651_inst_req_1;
      RPIPE_Block3_start_2593_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2596_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2599_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2602_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2605_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2608_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2611_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2614_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2617_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2620_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2633_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2645_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2648_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2651_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2594 <= data_out(223 downto 208);
      call1_2597 <= data_out(207 downto 192);
      call3_2600 <= data_out(191 downto 176);
      call5_2603 <= data_out(175 downto 160);
      call7_2606 <= data_out(159 downto 144);
      call9_2609 <= data_out(143 downto 128);
      call11_2612 <= data_out(127 downto 112);
      call13_2615 <= data_out(111 downto 96);
      call14_2618 <= data_out(95 downto 80);
      call15_2621 <= data_out(79 downto 64);
      call16_2634 <= data_out(63 downto 48);
      call18_2646 <= data_out(47 downto 32);
      call20_2649 <= data_out(31 downto 16);
      call22_2652 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2940_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2940_inst_req_0;
      WPIPE_Block3_done_2940_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2940_inst_req_1;
      WPIPE_Block3_done_2940_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2942_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_resp_35_inst_req_0 : boolean;
  signal RPIPE_timer_resp_35_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_35_inst_req_1 : boolean;
  signal WPIPE_timer_req_30_inst_req_0 : boolean;
  signal WPIPE_timer_req_30_inst_ack_0 : boolean;
  signal WPIPE_timer_req_30_inst_req_1 : boolean;
  signal WPIPE_timer_req_30_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_35_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_sample_start_
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/$entry
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_sample_start_
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Sample/req
      -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_30_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_35_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_sample_completed_
      -- CP-element group 1: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_update_start_
      -- CP-element group 1: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Sample/ack
      -- CP-element group 1: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Update/$entry
      -- CP-element group 1: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_30_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_30_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_update_completed_
      -- CP-element group 2: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Update/$exit
      -- CP-element group 2: 	 assign_stmt_33_to_assign_stmt_36/WPIPE_timer_req_30_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_30_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_sample_completed_
      -- CP-element group 3: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_update_start_
      -- CP-element group 3: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Sample/ra
      -- CP-element group 3: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Update/$entry
      -- CP-element group 3: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_35_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_35_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_update_completed_
      -- CP-element group 4: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Update/$exit
      -- CP-element group 4: 	 assign_stmt_33_to_assign_stmt_36/RPIPE_timer_resp_35_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_35_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_33_to_assign_stmt_36/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(2) & timer_CP_0_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_32_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_32_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_35_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_35_inst_req_0;
      RPIPE_timer_resp_35_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_35_inst_req_1;
      RPIPE_timer_resp_35_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_30_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_30_inst_req_0;
      WPIPE_timer_req_30_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_30_inst_req_1;
      WPIPE_timer_req_30_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_32_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    timer_req_pipe_read_data: out std_logic_vector(0 downto 0);
    timer_req_pipe_read_req : in std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : out std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data: in std_logic_vector(63 downto 0);
    timer_resp_pipe_write_req : in std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(10 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(69 downto 56),
      memory_space_2_sr_data => memory_space_2_sr_data(319 downto 256),
      memory_space_2_sr_tag => memory_space_2_sr_tag(94 downto 76),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(41 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(56 downto 38),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(191 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(2 downto 2),
      memory_space_2_sr_ack => memory_space_2_sr_ack(2 downto 2),
      memory_space_2_sr_addr => memory_space_2_sr_addr(41 downto 28),
      memory_space_2_sr_data => memory_space_2_sr_data(191 downto 128),
      memory_space_2_sr_tag => memory_space_2_sr_tag(56 downto 38),
      memory_space_2_sc_req => memory_space_2_sc_req(2 downto 2),
      memory_space_2_sc_ack => memory_space_2_sc_ack(2 downto 2),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 2),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(55 downto 42),
      memory_space_0_lr_tag => memory_space_0_lr_tag(75 downto 57),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(255 downto 192),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 3),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 3),
      memory_space_2_sr_addr => memory_space_2_sr_addr(55 downto 42),
      memory_space_2_sr_data => memory_space_2_sr_data(255 downto 192),
      memory_space_2_sr_tag => memory_space_2_sr_tag(75 downto 57),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 3),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 3),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 3),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 1),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(27 downto 14),
      memory_space_2_sr_data => memory_space_2_sr_data(127 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(37 downto 19),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
