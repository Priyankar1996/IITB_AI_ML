-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_728_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1011_inst_req_0 : boolean;
  signal type_cast_728_inst_req_1 : boolean;
  signal type_cast_728_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1064_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1348_inst_req_0 : boolean;
  signal type_cast_660_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1076_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1064_inst_req_1 : boolean;
  signal type_cast_575_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1064_inst_ack_1 : boolean;
  signal type_cast_611_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1073_inst_req_0 : boolean;
  signal type_cast_728_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1085_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1064_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 : boolean;
  signal type_cast_1056_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_req_1 : boolean;
  signal type_cast_575_inst_req_1 : boolean;
  signal type_cast_660_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1354_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal ptr_deref_619_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_ack_1 : boolean;
  signal type_cast_660_inst_ack_1 : boolean;
  signal type_cast_39_inst_req_0 : boolean;
  signal type_cast_39_inst_ack_0 : boolean;
  signal type_cast_39_inst_req_1 : boolean;
  signal ptr_deref_619_store_0_req_0 : boolean;
  signal type_cast_39_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 : boolean;
  signal type_cast_52_inst_req_0 : boolean;
  signal type_cast_52_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1070_inst_ack_0 : boolean;
  signal type_cast_52_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 : boolean;
  signal type_cast_575_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_ack_1 : boolean;
  signal type_cast_660_inst_req_1 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal addr_of_690_final_reg_ack_0 : boolean;
  signal type_cast_575_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1045_inst_ack_1 : boolean;
  signal type_cast_697_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1366_inst_req_1 : boolean;
  signal type_cast_77_inst_req_0 : boolean;
  signal type_cast_77_inst_ack_0 : boolean;
  signal type_cast_77_inst_req_1 : boolean;
  signal type_cast_77_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 : boolean;
  signal type_cast_710_inst_ack_1 : boolean;
  signal type_cast_697_inst_req_1 : boolean;
  signal type_cast_89_inst_req_0 : boolean;
  signal type_cast_89_inst_ack_0 : boolean;
  signal type_cast_89_inst_req_1 : boolean;
  signal type_cast_89_inst_ack_1 : boolean;
  signal addr_of_690_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1067_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 : boolean;
  signal type_cast_697_inst_ack_0 : boolean;
  signal type_cast_697_inst_req_0 : boolean;
  signal array_obj_ref_689_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1035_inst_req_1 : boolean;
  signal type_cast_102_inst_req_0 : boolean;
  signal type_cast_102_inst_ack_0 : boolean;
  signal type_cast_102_inst_req_1 : boolean;
  signal type_cast_102_inst_ack_1 : boolean;
  signal addr_of_690_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_ack_1 : boolean;
  signal addr_of_690_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 : boolean;
  signal type_cast_710_inst_req_1 : boolean;
  signal array_obj_ref_689_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_req_0 : boolean;
  signal type_cast_114_inst_req_0 : boolean;
  signal type_cast_114_inst_ack_0 : boolean;
  signal type_cast_114_inst_req_1 : boolean;
  signal type_cast_114_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1045_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_ack_1 : boolean;
  signal type_cast_127_inst_req_0 : boolean;
  signal type_cast_127_inst_ack_0 : boolean;
  signal type_cast_127_inst_req_1 : boolean;
  signal type_cast_127_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_ack_1 : boolean;
  signal if_stmt_633_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_1011_inst_req_1 : boolean;
  signal type_cast_340_inst_req_0 : boolean;
  signal type_cast_340_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1005_inst_req_0 : boolean;
  signal type_cast_340_inst_req_1 : boolean;
  signal type_cast_340_inst_ack_1 : boolean;
  signal type_cast_1306_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1014_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_349_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1014_inst_ack_1 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1067_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_req_0 : boolean;
  signal type_cast_152_inst_req_0 : boolean;
  signal type_cast_152_inst_ack_0 : boolean;
  signal type_cast_152_inst_req_1 : boolean;
  signal type_cast_152_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_req_1 : boolean;
  signal if_stmt_633_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 : boolean;
  signal type_cast_710_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1348_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_req_1 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_ack_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_1 : boolean;
  signal WPIPE_Block0_start_997_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 : boolean;
  signal array_obj_ref_689_index_offset_ack_0 : boolean;
  signal WPIPE_Block1_start_1020_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_req_1 : boolean;
  signal type_cast_177_inst_req_0 : boolean;
  signal type_cast_177_inst_ack_0 : boolean;
  signal type_cast_177_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_ack_0 : boolean;
  signal type_cast_177_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 : boolean;
  signal type_cast_557_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_0 : boolean;
  signal type_cast_189_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_1 : boolean;
  signal type_cast_189_inst_ack_1 : boolean;
  signal type_cast_557_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 : boolean;
  signal type_cast_710_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_607_inst_req_0 : boolean;
  signal type_cast_202_inst_req_0 : boolean;
  signal type_cast_202_inst_ack_0 : boolean;
  signal type_cast_202_inst_req_1 : boolean;
  signal type_cast_202_inst_ack_1 : boolean;
  signal type_cast_557_inst_ack_0 : boolean;
  signal type_cast_557_inst_req_0 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_req_1 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_0 : boolean;
  signal type_cast_215_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_1 : boolean;
  signal type_cast_215_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_ack_1 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal type_cast_521_inst_ack_1 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_ack_1 : boolean;
  signal type_cast_256_inst_req_0 : boolean;
  signal type_cast_256_inst_ack_0 : boolean;
  signal type_cast_521_inst_req_1 : boolean;
  signal type_cast_256_inst_req_1 : boolean;
  signal type_cast_256_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1082_inst_ack_1 : boolean;
  signal type_cast_260_inst_req_0 : boolean;
  signal type_cast_260_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_1 : boolean;
  signal type_cast_260_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_ack_0 : boolean;
  signal ptr_deref_619_store_0_ack_1 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal type_cast_264_inst_req_0 : boolean;
  signal type_cast_264_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1035_inst_ack_0 : boolean;
  signal type_cast_264_inst_req_1 : boolean;
  signal type_cast_264_inst_ack_1 : boolean;
  signal type_cast_1056_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_req_0 : boolean;
  signal ptr_deref_619_store_0_req_1 : boolean;
  signal type_cast_268_inst_req_0 : boolean;
  signal type_cast_268_inst_ack_0 : boolean;
  signal type_cast_521_inst_ack_0 : boolean;
  signal type_cast_268_inst_req_1 : boolean;
  signal type_cast_268_inst_ack_1 : boolean;
  signal if_stmt_633_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1011_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_286_inst_ack_1 : boolean;
  signal array_obj_ref_689_index_offset_req_0 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal type_cast_290_inst_req_0 : boolean;
  signal type_cast_290_inst_ack_0 : boolean;
  signal type_cast_290_inst_req_1 : boolean;
  signal type_cast_290_inst_ack_1 : boolean;
  signal type_cast_539_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_req_0 : boolean;
  signal WPIPE_Block0_start_997_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_ack_0 : boolean;
  signal type_cast_539_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_299_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_req_0 : boolean;
  signal type_cast_303_inst_req_0 : boolean;
  signal type_cast_611_inst_ack_1 : boolean;
  signal type_cast_303_inst_ack_0 : boolean;
  signal type_cast_303_inst_req_1 : boolean;
  signal type_cast_303_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_req_0 : boolean;
  signal type_cast_611_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_ack_0 : boolean;
  signal type_cast_539_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_311_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1038_inst_ack_0 : boolean;
  signal type_cast_315_inst_req_0 : boolean;
  signal type_cast_315_inst_ack_0 : boolean;
  signal type_cast_315_inst_req_1 : boolean;
  signal type_cast_315_inst_ack_1 : boolean;
  signal type_cast_539_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_req_1 : boolean;
  signal type_cast_611_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_324_inst_ack_1 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_req_1 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal type_cast_328_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1038_inst_ack_1 : boolean;
  signal type_cast_328_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1014_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1014_inst_ack_0 : boolean;
  signal type_cast_353_inst_req_0 : boolean;
  signal type_cast_353_inst_ack_0 : boolean;
  signal type_cast_353_inst_req_1 : boolean;
  signal type_cast_353_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_361_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1005_inst_ack_0 : boolean;
  signal type_cast_365_inst_req_0 : boolean;
  signal type_cast_365_inst_ack_0 : boolean;
  signal type_cast_365_inst_req_1 : boolean;
  signal type_cast_365_inst_ack_1 : boolean;
  signal type_cast_1056_inst_req_1 : boolean;
  signal type_cast_1043_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_374_inst_ack_1 : boolean;
  signal type_cast_378_inst_req_0 : boolean;
  signal type_cast_378_inst_ack_0 : boolean;
  signal type_cast_378_inst_req_1 : boolean;
  signal type_cast_378_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_386_inst_ack_1 : boolean;
  signal type_cast_1043_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1017_inst_req_0 : boolean;
  signal type_cast_390_inst_req_0 : boolean;
  signal type_cast_390_inst_ack_0 : boolean;
  signal type_cast_390_inst_req_1 : boolean;
  signal type_cast_390_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1017_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_399_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1070_inst_req_0 : boolean;
  signal type_cast_1306_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1079_inst_req_1 : boolean;
  signal type_cast_403_inst_req_0 : boolean;
  signal type_cast_403_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1020_inst_ack_1 : boolean;
  signal type_cast_403_inst_req_1 : boolean;
  signal type_cast_403_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1079_inst_ack_1 : boolean;
  signal if_stmt_417_branch_req_0 : boolean;
  signal if_stmt_417_branch_ack_1 : boolean;
  signal if_stmt_417_branch_ack_0 : boolean;
  signal if_stmt_432_branch_req_0 : boolean;
  signal if_stmt_432_branch_ack_1 : boolean;
  signal if_stmt_432_branch_ack_0 : boolean;
  signal type_cast_453_inst_req_0 : boolean;
  signal type_cast_453_inst_ack_0 : boolean;
  signal type_cast_453_inst_req_1 : boolean;
  signal type_cast_453_inst_ack_1 : boolean;
  signal array_obj_ref_482_index_offset_req_0 : boolean;
  signal array_obj_ref_482_index_offset_ack_0 : boolean;
  signal array_obj_ref_482_index_offset_req_1 : boolean;
  signal array_obj_ref_482_index_offset_ack_1 : boolean;
  signal addr_of_483_final_reg_req_0 : boolean;
  signal addr_of_483_final_reg_ack_0 : boolean;
  signal addr_of_483_final_reg_req_1 : boolean;
  signal addr_of_483_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_ack_1 : boolean;
  signal type_cast_490_inst_req_0 : boolean;
  signal type_cast_490_inst_ack_0 : boolean;
  signal type_cast_490_inst_req_1 : boolean;
  signal type_cast_490_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 : boolean;
  signal type_cast_503_inst_req_0 : boolean;
  signal type_cast_503_inst_ack_0 : boolean;
  signal type_cast_503_inst_req_1 : boolean;
  signal type_cast_503_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_ack_1 : boolean;
  signal type_cast_521_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1079_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1032_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1085_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_ack_0 : boolean;
  signal type_cast_746_inst_req_0 : boolean;
  signal type_cast_746_inst_ack_0 : boolean;
  signal type_cast_746_inst_req_1 : boolean;
  signal type_cast_746_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1366_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_req_0 : boolean;
  signal type_cast_764_inst_req_0 : boolean;
  signal type_cast_764_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_req_0 : boolean;
  signal type_cast_764_inst_req_1 : boolean;
  signal type_cast_764_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1366_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1061_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1061_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1348_inst_ack_0 : boolean;
  signal type_cast_782_inst_req_0 : boolean;
  signal type_cast_782_inst_ack_0 : boolean;
  signal type_cast_782_inst_req_1 : boolean;
  signal type_cast_782_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1008_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1076_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1061_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1008_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1061_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_req_1 : boolean;
  signal type_cast_800_inst_req_0 : boolean;
  signal type_cast_800_inst_ack_0 : boolean;
  signal type_cast_800_inst_req_1 : boolean;
  signal type_cast_800_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1029_inst_ack_0 : boolean;
  signal type_cast_476_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_814_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1008_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1091_inst_req_0 : boolean;
  signal type_cast_476_inst_req_1 : boolean;
  signal type_cast_818_inst_req_0 : boolean;
  signal type_cast_818_inst_ack_0 : boolean;
  signal type_cast_818_inst_req_1 : boolean;
  signal type_cast_818_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1058_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1058_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1017_inst_ack_1 : boolean;
  signal ptr_deref_826_store_0_req_0 : boolean;
  signal ptr_deref_826_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1045_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1001_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1017_inst_req_1 : boolean;
  signal ptr_deref_826_store_0_req_1 : boolean;
  signal WPIPE_Block1_start_1026_inst_ack_1 : boolean;
  signal ptr_deref_826_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_1026_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1045_inst_req_0 : boolean;
  signal if_stmt_840_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1001_inst_ack_0 : boolean;
  signal if_stmt_840_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_req_0 : boolean;
  signal if_stmt_840_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_req_0 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1008_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1070_inst_ack_1 : boolean;
  signal type_cast_855_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1058_inst_ack_0 : boolean;
  signal type_cast_855_inst_ack_0 : boolean;
  signal type_cast_855_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1058_inst_req_0 : boolean;
  signal type_cast_855_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1070_inst_req_1 : boolean;
  signal type_cast_859_inst_req_0 : boolean;
  signal type_cast_859_inst_ack_0 : boolean;
  signal ptr_deref_1272_load_0_ack_1 : boolean;
  signal type_cast_859_inst_req_1 : boolean;
  signal type_cast_859_inst_ack_1 : boolean;
  signal if_stmt_877_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1023_inst_ack_1 : boolean;
  signal type_cast_1043_inst_ack_1 : boolean;
  signal if_stmt_877_branch_ack_1 : boolean;
  signal if_stmt_877_branch_ack_0 : boolean;
  signal type_cast_1043_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_req_1 : boolean;
  signal type_cast_904_inst_req_0 : boolean;
  signal type_cast_904_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_1 : boolean;
  signal type_cast_904_inst_req_1 : boolean;
  signal type_cast_904_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1005_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1005_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1348_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1023_inst_req_0 : boolean;
  signal WPIPE_Block0_start_994_inst_req_1 : boolean;
  signal array_obj_ref_933_index_offset_req_0 : boolean;
  signal type_cast_1056_inst_ack_1 : boolean;
  signal array_obj_ref_933_index_offset_ack_0 : boolean;
  signal array_obj_ref_933_index_offset_req_1 : boolean;
  signal array_obj_ref_933_index_offset_ack_1 : boolean;
  signal type_cast_476_inst_ack_1 : boolean;
  signal type_cast_1306_inst_req_1 : boolean;
  signal addr_of_934_final_reg_req_0 : boolean;
  signal addr_of_934_final_reg_ack_0 : boolean;
  signal addr_of_934_final_reg_req_1 : boolean;
  signal addr_of_934_final_reg_ack_1 : boolean;
  signal phi_stmt_470_req_1 : boolean;
  signal ptr_deref_1272_load_0_req_0 : boolean;
  signal ptr_deref_1272_load_0_ack_0 : boolean;
  signal type_cast_1306_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1369_inst_req_0 : boolean;
  signal ptr_deref_937_store_0_req_0 : boolean;
  signal ptr_deref_937_store_0_ack_0 : boolean;
  signal ptr_deref_937_store_0_req_1 : boolean;
  signal ptr_deref_937_store_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1351_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1351_inst_ack_0 : boolean;
  signal if_stmt_952_branch_req_0 : boolean;
  signal if_stmt_952_branch_ack_1 : boolean;
  signal if_stmt_952_branch_ack_0 : boolean;
  signal call_stmt_963_call_req_0 : boolean;
  signal call_stmt_963_call_ack_0 : boolean;
  signal call_stmt_963_call_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1351_inst_req_1 : boolean;
  signal call_stmt_963_call_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1354_inst_ack_0 : boolean;
  signal type_cast_968_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1351_inst_ack_1 : boolean;
  signal type_cast_968_inst_ack_0 : boolean;
  signal type_cast_968_inst_req_1 : boolean;
  signal type_cast_968_inst_ack_1 : boolean;
  signal type_cast_476_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1369_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_1 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_973_inst_req_0 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_973_inst_req_1 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_976_inst_req_0 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_976_inst_req_1 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_979_inst_req_0 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_979_inst_req_1 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_982_inst_req_0 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_982_inst_req_1 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_985_inst_req_0 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_985_inst_req_1 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_req_0 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_988_inst_req_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_991_inst_req_0 : boolean;
  signal WPIPE_Block0_start_991_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_991_inst_req_1 : boolean;
  signal WPIPE_Block0_start_991_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_req_0 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_0 : boolean;
  signal type_cast_1099_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1366_inst_req_0 : boolean;
  signal type_cast_1099_inst_ack_0 : boolean;
  signal type_cast_1099_inst_req_1 : boolean;
  signal type_cast_1099_inst_ack_1 : boolean;
  signal type_cast_1346_inst_ack_1 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1101_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1101_inst_ack_0 : boolean;
  signal ptr_deref_1272_load_0_req_1 : boolean;
  signal WPIPE_Block2_start_1101_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1101_inst_ack_1 : boolean;
  signal type_cast_1112_inst_req_0 : boolean;
  signal type_cast_1112_inst_ack_0 : boolean;
  signal type_cast_1112_inst_req_1 : boolean;
  signal type_cast_1112_inst_ack_1 : boolean;
  signal if_stmt_1383_branch_ack_0 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1114_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1114_inst_ack_0 : boolean;
  signal type_cast_1296_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1114_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1114_inst_ack_1 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1117_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1363_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1117_inst_ack_0 : boolean;
  signal type_cast_1296_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1117_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1363_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1117_inst_ack_1 : boolean;
  signal if_stmt_1383_branch_ack_1 : boolean;
  signal WPIPE_Block2_start_1120_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1120_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1120_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1120_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1123_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1363_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1363_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1126_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1126_inst_ack_0 : boolean;
  signal type_cast_1296_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1126_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1126_inst_ack_1 : boolean;
  signal if_stmt_1383_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1129_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1129_inst_ack_0 : boolean;
  signal type_cast_1296_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1129_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1129_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1132_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1132_inst_ack_1 : boolean;
  signal type_cast_1336_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1360_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1135_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1360_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_ack_1 : boolean;
  signal type_cast_1336_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1138_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1138_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1141_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1360_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1141_inst_ack_1 : boolean;
  signal phi_stmt_470_req_0 : boolean;
  signal WPIPE_Block3_start_1144_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1360_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1144_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1144_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1144_inst_ack_1 : boolean;
  signal phi_stmt_677_ack_0 : boolean;
  signal type_cast_1336_inst_ack_0 : boolean;
  signal type_cast_1336_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1147_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1147_inst_ack_0 : boolean;
  signal type_cast_1286_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_ack_1 : boolean;
  signal type_cast_1286_inst_req_1 : boolean;
  signal phi_stmt_677_req_1 : boolean;
  signal type_cast_683_inst_ack_1 : boolean;
  signal type_cast_683_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1150_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1150_inst_ack_1 : boolean;
  signal type_cast_683_inst_ack_0 : boolean;
  signal type_cast_1155_inst_req_0 : boolean;
  signal type_cast_1155_inst_ack_0 : boolean;
  signal phi_stmt_470_ack_0 : boolean;
  signal type_cast_1155_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1357_inst_ack_1 : boolean;
  signal type_cast_1155_inst_ack_1 : boolean;
  signal type_cast_1286_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1369_inst_ack_1 : boolean;
  signal type_cast_1286_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1369_inst_req_1 : boolean;
  signal type_cast_1326_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1157_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1357_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1157_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1157_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1157_inst_ack_1 : boolean;
  signal type_cast_683_inst_req_0 : boolean;
  signal type_cast_1326_inst_req_1 : boolean;
  signal type_cast_1326_inst_ack_0 : boolean;
  signal type_cast_1168_inst_req_0 : boolean;
  signal type_cast_1168_inst_ack_0 : boolean;
  signal type_cast_1168_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1357_inst_ack_0 : boolean;
  signal type_cast_1168_inst_ack_1 : boolean;
  signal type_cast_1326_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1170_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1357_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1170_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1170_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1170_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1173_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1173_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1173_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1173_inst_ack_1 : boolean;
  signal type_cast_1276_inst_ack_1 : boolean;
  signal type_cast_1316_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1176_inst_ack_0 : boolean;
  signal type_cast_1276_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_ack_1 : boolean;
  signal type_cast_1316_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1179_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1179_inst_ack_1 : boolean;
  signal type_cast_1276_inst_ack_0 : boolean;
  signal phi_stmt_677_req_0 : boolean;
  signal type_cast_1316_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1183_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1354_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1183_inst_ack_0 : boolean;
  signal type_cast_1276_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1183_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1354_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1183_inst_ack_1 : boolean;
  signal type_cast_1316_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1186_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1186_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1186_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1186_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1189_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1189_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1189_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1189_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1192_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1192_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1192_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1192_inst_ack_1 : boolean;
  signal call_stmt_1196_call_req_0 : boolean;
  signal call_stmt_1196_call_ack_0 : boolean;
  signal call_stmt_1196_call_req_1 : boolean;
  signal call_stmt_1196_call_ack_1 : boolean;
  signal type_cast_1200_inst_req_0 : boolean;
  signal type_cast_1200_inst_ack_0 : boolean;
  signal type_cast_1200_inst_req_1 : boolean;
  signal type_cast_1200_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1207_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1207_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1207_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1207_inst_ack_1 : boolean;
  signal if_stmt_1211_branch_req_0 : boolean;
  signal if_stmt_1211_branch_ack_1 : boolean;
  signal if_stmt_1211_branch_ack_0 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal array_obj_ref_1267_index_offset_req_0 : boolean;
  signal array_obj_ref_1267_index_offset_ack_0 : boolean;
  signal array_obj_ref_1267_index_offset_req_1 : boolean;
  signal array_obj_ref_1267_index_offset_ack_1 : boolean;
  signal addr_of_1268_final_reg_req_0 : boolean;
  signal addr_of_1268_final_reg_ack_0 : boolean;
  signal addr_of_1268_final_reg_req_1 : boolean;
  signal addr_of_1268_final_reg_ack_1 : boolean;
  signal phi_stmt_921_req_1 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_1 : boolean;
  signal type_cast_924_inst_ack_1 : boolean;
  signal phi_stmt_921_req_0 : boolean;
  signal phi_stmt_921_ack_0 : boolean;
  signal phi_stmt_1255_req_0 : boolean;
  signal type_cast_1261_inst_req_0 : boolean;
  signal type_cast_1261_inst_ack_0 : boolean;
  signal type_cast_1261_inst_req_1 : boolean;
  signal type_cast_1261_inst_ack_1 : boolean;
  signal phi_stmt_1255_req_1 : boolean;
  signal phi_stmt_1255_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(459 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(459);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_33/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/branch_block_stmt_33__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/cr
      -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_39_inst_req_1); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_52_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_64_inst_req_1); -- 
    cr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_77_inst_req_1); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_89_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_102_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_114_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_127_inst_req_1); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_340_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_139_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_152_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_164_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_177_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_189_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_202_inst_req_1); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_215_inst_req_1); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_219_inst_req_1); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_256_inst_req_1); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_260_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_264_inst_req_1); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_268_inst_req_1); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_290_inst_req_1); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_303_inst_req_1); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_315_inst_req_1); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_328_inst_req_1); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_353_inst_req_1); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_365_inst_req_1); -- 
    cr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_378_inst_req_1); -- 
    cr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_390_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_403_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/rr
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_39_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Sample/ra
      -- 
    ra_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_39_Update/ca
      -- 
    ca_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_update_start_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/cr
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_48_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/rr
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_52_inst_req_0); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Sample/ra
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_52_Update/ca
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_update_start_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/cr
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_60_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/rr
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_64_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_64_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_update_start_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_73_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_77_inst_req_0); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Sample/ra
      -- 
    ra_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_77_Update/ca
      -- 
    ca_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_update_start_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_85_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_0); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_89_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_89_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_update_start_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_98_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_102_inst_req_0); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_102_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_update_start_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_110_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_0); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_114_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_114_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_update_start_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_123_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/$entry
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_127_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_127_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_update_start_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Sample/$exit
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_135_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_139_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_139_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_update_start_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_148_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_152_inst_req_0); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_152_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_update_start_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_160_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_164_inst_req_0); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_164_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_update_start_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_173_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_177_inst_req_0); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_177_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_update_start_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_185_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_189_inst_req_0); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_189_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_update_start_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_198_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_202_inst_req_0); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_286_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_202_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/rr
      -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_211_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Sample/ra
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_211_Update/ca
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/rr
      -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_215_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_215_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	24 
    -- CP-element group 63: 	20 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/rr
      -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_219_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(24) & convTranspose_CP_39_elements(20);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Sample/ra
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_219_Update/ca
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/rr
      -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_256_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Sample/ra
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_256_Update/ca
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/rr
      -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_260_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Sample/ra
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_260_Update/ca
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/rr
      -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_264_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(44) & convTranspose_CP_39_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_264_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/rr
      -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_268_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Sample/ra
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_268_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_268_Update/ca
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_268_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_update_start_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/cr
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_286_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_286_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_286_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/rr
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_286_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_290_inst_req_0); -- 
    rr_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_299_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Sample/ra
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_290_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_290_Update/ca
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_290_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_update_start_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/cr
      -- 
    ra_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_299_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_299_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_299_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/rr
      -- 
    ca_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_299_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_303_inst_req_0); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_311_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Sample/ra
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_303_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_303_Update/ca
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_303_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_update_start_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/cr
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_311_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_311_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_311_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/rr
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_311_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_315_inst_req_0); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_324_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Sample/ra
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_315_Update/ca
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_update_start_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/cr
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_324_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_324_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_324_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/rr
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_324_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_328_inst_req_0); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Sample/ra
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_328_Update/ca
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_328_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_update_start_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/cr
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_336_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_336_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_sample_start_
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_336_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_340_inst_req_0); -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_349_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_sample_completed_
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_340_update_completed_
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_update_start_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/cr
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_349_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_349_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_349_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/rr
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_349_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_353_inst_req_0); -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_361_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Sample/ra
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_353_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_353_Update/ca
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_353_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_update_start_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/cr
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_361_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_361_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_361_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/rr
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_361_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_365_inst_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_374_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Sample/ra
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_365_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_365_Update/ca
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_365_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_update_start_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/cr
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_374_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_374_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_374_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/rr
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_374_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_378_inst_req_0); -- 
    rr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_386_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Sample/ra
      -- 
    ra_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_378_Update/ca
      -- 
    ca_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_378_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_update_start_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/cr
      -- 
    ra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_386_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_386_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_386_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/rr
      -- 
    ca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_386_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_390_inst_req_0); -- 
    rr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_399_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Sample/ra
      -- 
    ra_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_390_Update/ca
      -- 
    ca_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_update_start_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/cr
      -- 
    ra_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_399_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_399_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/RPIPE_ConvTranspose_input_pipe_399_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/rr
      -- 
    ca_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_399_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_403_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Sample/ra
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/type_cast_403_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416__exit__
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417__entry__
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_416/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_33/R_cmp451_418_place
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_417_else_link/$entry
      -- 
    branch_req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_417_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(117) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438__exit__
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467__entry__
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_417_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_417_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph453
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_update_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph453_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph453_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_438_PhiAck/dummy
      -- 
    if_choice_transition_908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_417_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_453_inst_req_0); -- 
    cr_952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_453_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	432 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_417_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_417_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond190x_xpreheader
      -- 
    else_choice_transition_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_417_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	432 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639__exit__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674__entry__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_update_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_432_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_432_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_bbx_xnph449
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiAck/dummy
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_639_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_bbx_xnph449_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_bbx_xnph449_PhiReq/$entry
      -- 
    if_choice_transition_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_432_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_660_inst_req_0); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_660_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	432 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	445 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_432_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_432_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- 
    else_choice_transition_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_432_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Sample/ra
      -- 
    ra_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	433 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467__exit__
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_444_to_assign_stmt_467/type_cast_453_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/phi_stmt_470/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/$entry
      -- 
    ca_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_453_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	438 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/ack
      -- 
    ack_982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_482_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	438 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/req
      -- 
    ack_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_482_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_483_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_request/ack
      -- 
    ack_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_483_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	438 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/ack
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_483_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	438 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_update_start_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/cr
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_486_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_486_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/rr
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_486_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_490_inst_req_0); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Sample/ra
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	438 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/ca
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_update_start_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/cr
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_499_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/rr
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_503_inst_req_0); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_517_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Sample/ra
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	438 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/ca
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_update_start_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/cr
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_517_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_517_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	141 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_517_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/rr
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_517_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_521_inst_req_0); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_535_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Sample/$exit
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_521_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	438 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_update_completed_
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_521_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_update_start_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_sample_completed_
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_535_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_535_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_535_update_completed_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_535_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_539_inst_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_553_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Sample/$exit
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	438 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/$exit
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_update_start_
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_sample_completed_
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_553_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_553_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_553_update_completed_
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_553_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_557_inst_req_0); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_571_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_sample_completed_
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_557_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	438 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_update_completed_
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_557_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_update_start_
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_sample_completed_
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_571_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_571_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_571_update_completed_
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_571_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_575_inst_req_0); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_589_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Sample/$exit
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_575_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	438 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_update_completed_
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_575_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_update_start_
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_589_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_589_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_589_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/$entry
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_589_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_593_inst_req_0); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_607_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_sample_completed_
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	438 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_update_completed_
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_update_start_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_sample_completed_
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_607_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_607_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_607_update_completed_
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_607_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_611_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Sample/ra
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	438 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/$exit
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/ptr_deref_619_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_sample_start_
      -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_619_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(156) & convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_sample_completed_
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	438 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/$exit
      -- 
    ca_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632__exit__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633__entry__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/R_exitcond3_634_place
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_633_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/$exit
      -- 
    branch_req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_633_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	432 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423__exit__
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_633_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_633_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_423_PhiReqMerge
      -- 
    if_choice_transition_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_633_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	434 
    -- CP-element group 166: 	435 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_633_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_633_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/cr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_633_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    rr_3296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_476_inst_req_0); -- 
    cr_3301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_476_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_sample_completed_
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	439 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674__exit__
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_645_to_assign_stmt_674/type_cast_660_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/phi_stmt_677/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$entry
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	444 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_sample_complete
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/$exit
      -- 
    ack_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_689_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	444 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_sample_start_
      -- 
    ack_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_689_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_690_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_sample_completed_
      -- 
    ack_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_690_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	444 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_word_addrgen/root_register_ack
      -- 
    ack_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_690_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	444 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_update_start_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/$exit
      -- 
    ra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_693_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_693_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_update_completed_
      -- 
    ca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_693_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_697_inst_req_0); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_706_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_sample_completed_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	444 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/$exit
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_update_start_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Sample/$exit
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_706_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_706_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_706_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/$entry
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_706_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_710_inst_req_0); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_724_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Sample/$exit
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_710_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	444 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_update_completed_
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_710_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_update_start_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/cr
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_724_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_724_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_724_Update/$exit
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_724_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_742_inst_req_0); -- 
    rr_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_728_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_sample_completed_
      -- 
    ra_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	444 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_update_completed_
      -- 
    ca_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_update_start_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/cr
      -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_742_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_742_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_742_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/rr
      -- 
    ca_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_742_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_746_inst_req_0); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Sample/ra
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_746_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	444 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/ca
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_746_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_update_start_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/cr
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_760_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/rr
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_764_inst_req_0); -- 
    rr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Sample/ra
      -- 
    ra_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	444 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/ca
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_update_start_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/cr
      -- 
    ra_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_778_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/rr
      -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_782_inst_req_0); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Sample/ra
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	444 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/ca
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_update_start_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/cr
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_796_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/rr
      -- 
    ca_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_800_inst_req_0); -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_814_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Sample/ra
      -- 
    ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	444 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/ca
      -- 
    ca_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_update_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/cr
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_814_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_814_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_814_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/rr
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_814_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_818_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Sample/ra
      -- 
    ra_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	444 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/ca
      -- 
    ca_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/ptr_deref_826_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/rr
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_826_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204) & convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Sample/word_access_start/word_0/ra
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_826_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	444 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/ca
      -- 
    ca_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_826_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839__exit__
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840__entry__
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_33/R_exitcond2_841_place
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_840_else_link/$entry
      -- 
    branch_req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_840_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(207) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	445 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846__exit__
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_840_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_840_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_846_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_840_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	440 
    -- CP-element group 210: 	441 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_840_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_840_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- 
    else_choice_transition_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_840_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    cr_3355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_683_inst_req_1); -- 
    rr_3350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_683_inst_req_0); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	445 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/ra
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	445 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/ca
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	445 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	445 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/ca
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	445 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/ra
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	445 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/ca
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876__exit__
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877__entry__
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_33/R_cmp264443_878_place
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_877_else_link/$entry
      -- 
    branch_req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_877_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883__exit__
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918__entry__
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_877_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_877_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend250_bbx_xnph445
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_update_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend250_bbx_xnph445_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend250_bbx_xnph445_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_883_PhiAck/dummy
      -- 
    if_choice_transition_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_877_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_904_inst_req_0); -- 
    cr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_904_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	452 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_877_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_877_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_877_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Sample/ra
      -- 
    ra_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_904_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	446 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918__exit__
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_889_to_assign_stmt_918/type_cast_904_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/phi_stmt_921/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$entry
      -- 
    ca_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_904_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	451 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/ack
      -- 
    ack_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_933_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	451 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/req
      -- 
    ack_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_933_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_934_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_request/ack
      -- 
    ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_934_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	451 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/ptr_deref_937_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/rr
      -- 
    ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_934_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_937_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Sample/word_access_start/word_0/ra
      -- 
    ra_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_937_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	451 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_937_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951__exit__
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952__entry__
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_33/R_exitcond_953_place
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_952_else_link/$entry
      -- 
    branch_req_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_952_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	452 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958__exit__
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_952_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_952_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_958_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_952_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	447 
    -- CP-element group 230: 	448 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_952_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_952_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_952_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_3427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_924_inst_req_0); -- 
    cr_3432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_924_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	452 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Sample/cra
      -- 
    cra_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_963_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	452 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Sample/rr
      -- 
    cca_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_963_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_968_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Sample/ra
      -- 
    ra_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	452 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	373 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Update/ca
      -- 
    ca_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	452 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_update_start_
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_970_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/req
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_973_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_update_start_
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/req
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_973_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/req
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_976_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_update_start_
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_976_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_979_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_update_start_
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_979_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/req
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_982_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_update_start_
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/req
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_982_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/req
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_985_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_update_start_
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/req
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_985_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/req
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_988_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_update_start_
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/req
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_988_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/req
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_991_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_991_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_991_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_991_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_994_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/req
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_update_start_
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/ack
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_994_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_994_update_completed_
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_997_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_update_start_
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/req
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/$exit
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_997_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_997_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/req
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_997_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_1001_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_update_start_
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/req
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/ack
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1001_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_1001_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/$exit
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1001_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_1005_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_update_start_
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/req
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1005_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_1005_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/ack
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1005_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block0_start_1008_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/req
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_update_start_
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_sample_completed_
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1008_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block0_start_1008_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1008_update_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1008_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block0_start_1011_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/req
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_update_start_
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_sample_completed_
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1011_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block0_start_1011_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_1011_update_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1011_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	452 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/req
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_update_start_
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/ack
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1014_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_1014_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/req
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1014_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_1017_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_update_start_
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/req
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1017_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_1017_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/ack
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1017_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1020_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/req
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1020_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1020_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_sample_start_
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1020_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1023_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/req
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_update_start_
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_sample_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1023_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1023_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1023_update_completed_
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1023_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1026_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/req
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_update_start_
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_sample_completed_
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1026_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1026_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1026_update_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1026_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1029_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/req
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_update_start_
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_sample_completed_
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1029_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1029_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1029_update_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1029_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1032_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/req
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_update_start_
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_sample_completed_
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1032_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1032_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1032_update_completed_
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1032_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1035_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/req
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_update_start_
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/ack
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1035_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1035_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/req
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1035_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1038_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_update_start_
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/req
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1038_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1038_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/ack
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1038_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	452 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Sample/ra
      -- 
    ra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1043_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	452 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Update/$exit
      -- 
    ca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1043_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_sample_start_
      -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block1_start_1045_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(280) & convTranspose_CP_39_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Update/req
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_update_start_
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_sample_completed_
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1045_inst_ack_0, ack => convTranspose_CP_39_elements(284)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block1_start_1045_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Update/ack
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1045_update_completed_
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1045_inst_ack_1, ack => convTranspose_CP_39_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	452 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Sample/ra
      -- 
    ra_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_0, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	452 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Update/ca
      -- 
    ca_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_1, ack => convTranspose_CP_39_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_sample_start_
      -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block1_start_1058_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(285) & convTranspose_CP_39_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/req
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_update_start_
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_sample_completed_
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1058_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block1_start_1058_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1058_update_completed_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1058_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block1_start_1061_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/req
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_update_start_
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_sample_completed_
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1061_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block1_start_1061_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1061_update_completed_
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1061_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block1_start_1064_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/req
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_update_start_
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_sample_completed_
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1064_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block1_start_1064_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1064_update_completed_
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1064_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block1_start_1067_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/req
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1067_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block1_start_1067_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1067_update_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1067_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	452 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_update_start_
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/req
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/$entry
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1070_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1070_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/$exit
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1070_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1073_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/req
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_update_start_
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_sample_completed_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1073_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1073_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1073_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/$entry
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1073_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1076_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/req
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/$exit
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1076_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1076_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/$entry
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1076_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1079_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/req
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_sample_completed_
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1079_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1079_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1079_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_sample_start_
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1079_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1082_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/req
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_update_start_
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_sample_completed_
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1082_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1082_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1082_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_sample_start_
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1082_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block2_start_1085_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/req
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_update_start_
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_sample_completed_
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1085_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block2_start_1085_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1085_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_sample_start_
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1085_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block2_start_1088_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_update_start_
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/req
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1088_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block2_start_1088_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/$exit
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1088_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block2_start_1091_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/req
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_update_start_
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/$exit
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1091_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block2_start_1091_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/req
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/ack
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1091_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block2_start_1094_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_update_start_
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/req
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/ack
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1094_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block2_start_1094_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/$exit
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1094_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	452 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Sample/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1099_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	452 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Update/ca
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1099_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Sample/req
      -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block2_start_1101_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(314) & convTranspose_CP_39_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_update_start_
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1101_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block2_start_1101_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1101_Update/ack
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1101_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	452 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	452 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Update/ca
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/req
      -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block2_start_1114_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_update_start_
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1114_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block2_start_1114_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1114_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block2_start_1117_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_update_start_
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1117_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block2_start_1117_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1117_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block2_start_1120_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_update_start_
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1120_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block2_start_1120_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1120_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block2_start_1123_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_update_start_
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1123_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block2_start_1123_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/ack
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1123_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	452 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_update_start_
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1126_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => WPIPE_Block3_start_1126_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1126_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(332), ack => WPIPE_Block3_start_1129_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_update_start_
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1129_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_Block3_start_1129_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1129_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_Block3_start_1132_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_update_start_
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1132_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => WPIPE_Block3_start_1132_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1132_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_Block3_start_1135_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_update_start_
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1135_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_Block3_start_1135_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1135_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(338), ack => WPIPE_Block3_start_1138_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_update_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1138_inst_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_Block3_start_1138_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1138_inst_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_Block3_start_1141_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_update_start_
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1141_inst_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => WPIPE_Block3_start_1141_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1141_inst_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_Block3_start_1144_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_update_start_
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1144_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_Block3_start_1144_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1144_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_Block3_start_1147_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_update_start_
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1147_inst_ack_0, ack => convTranspose_CP_39_elements(345)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_Block3_start_1147_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1147_inst_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_Block3_start_1150_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_update_start_
      -- CP-element group 347: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1150_inst_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => WPIPE_Block3_start_1150_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/ack
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1150_inst_ack_1, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	452 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Sample/ra
      -- 
    ra_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1155_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	452 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Update/ca
      -- 
    ca_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1155_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Sample/req
      -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_Block3_start_1157_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(348) & convTranspose_CP_39_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_update_start_
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Update/req
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1157_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block3_start_1157_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1157_Update/ack
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1157_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	452 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Sample/ra
      -- 
    ra_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	452 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Update/ca
      -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/req
      -- 
    req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(356), ack => WPIPE_Block3_start_1170_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(353) & convTranspose_CP_39_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_update_start_
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/req
      -- 
    ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1170_inst_ack_0, ack => convTranspose_CP_39_elements(357)); -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_Block3_start_1170_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1170_inst_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    req_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_Block3_start_1173_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_update_start_
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/req
      -- 
    ack_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1173_inst_ack_0, ack => convTranspose_CP_39_elements(359)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block3_start_1173_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1173_inst_ack_1, ack => convTranspose_CP_39_elements(360)); -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block3_start_1176_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_update_start_
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/req
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1176_inst_ack_0, ack => convTranspose_CP_39_elements(361)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_Block3_start_1176_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1176_inst_ack_1, ack => convTranspose_CP_39_elements(362)); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block3_start_1179_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_update_start_
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/req
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1179_inst_ack_0, ack => convTranspose_CP_39_elements(363)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block3_start_1179_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/ack
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1179_inst_ack_1, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	452 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_update_start_
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/cr
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1183_inst_ack_0, ack => convTranspose_CP_39_elements(365)); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => RPIPE_Block0_done_1183_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/ca
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1183_inst_ack_1, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	452 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_update_start_
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/cr
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1186_inst_ack_0, ack => convTranspose_CP_39_elements(367)); -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => RPIPE_Block1_done_1186_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/ca
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1186_inst_ack_1, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	452 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_update_start_
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/cr
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1189_inst_ack_0, ack => convTranspose_CP_39_elements(369)); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => RPIPE_Block2_done_1189_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/ca
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1189_inst_ack_1, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	452 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_update_start_
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/cr
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1192_inst_ack_0, ack => convTranspose_CP_39_elements(371)); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => RPIPE_Block3_done_1192_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1192_inst_ack_1, ack => convTranspose_CP_39_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	234 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: 	330 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	377 
    -- CP-element group 373:  members (13) 
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193__exit__
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209__entry__
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/$exit
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_update_start_
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Update/cr
      -- 
    crr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1196_call_req_0); -- 
    ccr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1196_call_req_1); -- 
    cr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1200_inst_req_1); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(234) & convTranspose_CP_39_elements(262) & convTranspose_CP_39_elements(296) & convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(364) & convTranspose_CP_39_elements(366) & convTranspose_CP_39_elements(368) & convTranspose_CP_39_elements(370) & convTranspose_CP_39_elements(372);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Sample/cra
      -- 
    cra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1196_call_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/call_stmt_1196_Update/cca
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Sample/rr
      -- 
    cca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1196_call_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    rr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => type_cast_1200_inst_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Sample/ra
      -- 
    ra_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/type_cast_1200_Update/ca
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Sample/req
      -- 
    ca_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    req_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => WPIPE_elapsed_time_pipe_1207_inst_req_0); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_update_start_
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Update/req
      -- 
    ack_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1207_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    req_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => WPIPE_elapsed_time_pipe_1207_inst_req_1); -- 
    -- CP-element group 379:  branch  transition  place  input  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (13) 
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209__exit__
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211__entry__
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/call_stmt_1196_to_assign_stmt_1209/WPIPE_elapsed_time_pipe_1207_Update/ack
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211_dead_link/$entry
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211_eval_test/$entry
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211_eval_test/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211_eval_test/branch_req
      -- CP-element group 379: 	 branch_block_stmt_33/R_cmp264443_1212_place
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211_if_link/$entry
      -- CP-element group 379: 	 branch_block_stmt_33/if_stmt_1211_else_link/$entry
      -- 
    ack_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1207_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    branch_req_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => if_stmt_1211_branch_req_0); -- 
    -- CP-element group 380:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: 	383 
    -- CP-element group 380:  members (18) 
      -- CP-element group 380: 	 branch_block_stmt_33/merge_stmt_1217__exit__
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252__entry__
      -- CP-element group 380: 	 branch_block_stmt_33/if_stmt_1211_if_link/$exit
      -- CP-element group 380: 	 branch_block_stmt_33/if_stmt_1211_if_link/if_choice_transition
      -- CP-element group 380: 	 branch_block_stmt_33/forx_xend273_bbx_xnph
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_update_start_
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Sample/rr
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Update/cr
      -- CP-element group 380: 	 branch_block_stmt_33/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 380: 	 branch_block_stmt_33/merge_stmt_1217_PhiReqMerge
      -- CP-element group 380: 	 branch_block_stmt_33/merge_stmt_1217_PhiAck/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/merge_stmt_1217_PhiAck/$exit
      -- CP-element group 380: 	 branch_block_stmt_33/merge_stmt_1217_PhiAck/dummy
      -- 
    if_choice_transition_2866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1211_branch_ack_1, ack => convTranspose_CP_39_elements(380)); -- 
    rr_2883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => type_cast_1238_inst_req_0); -- 
    cr_2888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => type_cast_1238_inst_req_1); -- 
    -- CP-element group 381:  transition  place  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	459 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 branch_block_stmt_33/if_stmt_1211_else_link/$exit
      -- CP-element group 381: 	 branch_block_stmt_33/if_stmt_1211_else_link/else_choice_transition
      -- CP-element group 381: 	 branch_block_stmt_33/forx_xend273_forx_xend438
      -- CP-element group 381: 	 branch_block_stmt_33/forx_xend273_forx_xend438_PhiReq/$entry
      -- CP-element group 381: 	 branch_block_stmt_33/forx_xend273_forx_xend438_PhiReq/$exit
      -- 
    else_choice_transition_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1211_branch_ack_0, ack => convTranspose_CP_39_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Sample/ra
      -- 
    ra_2884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  transition  place  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	380 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	453 
    -- CP-element group 383:  members (9) 
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252__exit__
      -- CP-element group 383: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/$exit
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1223_to_assign_stmt_1252/type_cast_1238_Update/ca
      -- CP-element group 383: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/$entry
      -- CP-element group 383: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/phi_stmt_1255/$entry
      -- CP-element group 383: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/$entry
      -- 
    ca_2889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	458 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	429 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_sample_complete
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Sample/ack
      -- 
    ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1267_index_offset_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    -- CP-element group 385:  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	458 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (11) 
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_root_address_calculated
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_offset_calculated
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Update/ack
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_base_plus_offset/$entry
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_base_plus_offset/$exit
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_base_plus_offset/sum_rename_req
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_base_plus_offset/sum_rename_ack
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_request/$entry
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_request/req
      -- 
    ack_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1267_index_offset_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    req_2932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(385), ack => addr_of_1268_final_reg_req_0); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_request/$exit
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_request/ack
      -- 
    ack_2933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1268_final_reg_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    -- CP-element group 387:  join  fork  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	458 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (24) 
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/word_access_start/word_0/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/word_access_start/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/word_access_start/word_0/rr
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_complete/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_complete/ack
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_address_calculated
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_word_address_calculated
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_root_address_calculated
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_address_resized
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_addr_resize/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_addr_resize/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_addr_resize/base_resize_req
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_addr_resize/base_resize_ack
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_plus_offset/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_plus_offset/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_plus_offset/sum_rename_req
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_base_plus_offset/sum_rename_ack
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_word_addrgen/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_word_addrgen/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_word_addrgen/root_register_req
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_word_addrgen/root_register_ack
      -- 
    ack_2938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1268_final_reg_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    rr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(387), ack => ptr_deref_1272_load_0_req_0); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (5) 
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/word_access_start/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/word_access_start/word_0/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Sample/word_access_start/word_0/ra
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_sample_completed_
      -- 
    ra_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1272_load_0_ack_0, ack => convTranspose_CP_39_elements(388)); -- 
    -- CP-element group 389:  fork  transition  input  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	458 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	404 
    -- CP-element group 389: 	390 
    -- CP-element group 389: 	392 
    -- CP-element group 389: 	394 
    -- CP-element group 389: 	396 
    -- CP-element group 389: 	398 
    -- CP-element group 389: 	400 
    -- CP-element group 389: 	402 
    -- CP-element group 389:  members (33) 
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/ptr_deref_1272_Merge/$exit
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/word_access_complete/word_0/ca
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/ptr_deref_1272_Merge/merge_req
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/ptr_deref_1272_Merge/merge_ack
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/ptr_deref_1272_Merge/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/word_access_complete/word_0/$exit
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/word_access_complete/$exit
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Sample/rr
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_update_completed_
      -- 
    ca_2983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1272_load_0_ack_1, ack => convTranspose_CP_39_elements(389)); -- 
    rr_3094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1346_inst_req_0); -- 
    rr_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1276_inst_req_0); -- 
    rr_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1286_inst_req_0); -- 
    rr_3024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1296_inst_req_0); -- 
    rr_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1306_inst_req_0); -- 
    rr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1316_inst_req_0); -- 
    rr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1326_inst_req_0); -- 
    rr_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => type_cast_1336_inst_req_0); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Sample/ra
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Sample/$exit
      -- 
    ra_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	458 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	426 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Update/ca
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Update/$exit
      -- 
    ca_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	389 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Sample/ra
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_sample_completed_
      -- 
    ra_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	458 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	423 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Update/ca
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_update_completed_
      -- 
    ca_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	389 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Sample/ra
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_sample_completed_
      -- 
    ra_3025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1296_inst_ack_0, ack => convTranspose_CP_39_elements(394)); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	458 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	420 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Update/ca
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_update_completed_
      -- 
    ca_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1296_inst_ack_1, ack => convTranspose_CP_39_elements(395)); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	389 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Sample/ra
      -- CP-element group 396: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_sample_completed_
      -- CP-element group 396: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Sample/$exit
      -- 
    ra_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1306_inst_ack_0, ack => convTranspose_CP_39_elements(396)); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	458 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	417 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_update_completed_
      -- CP-element group 397: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Update/ca
      -- 
    ca_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1306_inst_ack_1, ack => convTranspose_CP_39_elements(397)); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	389 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Sample/ra
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Sample/$exit
      -- 
    ra_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_0, ack => convTranspose_CP_39_elements(398)); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	458 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	414 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Update/ca
      -- CP-element group 399: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Update/$exit
      -- 
    ca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_1, ack => convTranspose_CP_39_elements(399)); -- 
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	389 
    -- CP-element group 400: successors 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Sample/ra
      -- CP-element group 400: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_sample_completed_
      -- 
    ra_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1326_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	458 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	411 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Update/ca
      -- CP-element group 401: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_update_completed_
      -- 
    ca_3072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1326_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	389 
    -- CP-element group 402: successors 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Sample/ra
      -- CP-element group 402: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_sample_completed_
      -- 
    ra_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_0, ack => convTranspose_CP_39_elements(402)); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	458 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	408 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Update/ca
      -- CP-element group 403: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Update/$exit
      -- CP-element group 403: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_update_completed_
      -- 
    ca_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_1, ack => convTranspose_CP_39_elements(403)); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	389 
    -- CP-element group 404: successors 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Sample/ra
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_sample_completed_
      -- 
    ra_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => convTranspose_CP_39_elements(404)); -- 
    -- CP-element group 405:  transition  input  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	458 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (6) 
      -- CP-element group 405: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Sample/req
      -- CP-element group 405: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_sample_start_
      -- CP-element group 405: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Update/ca
      -- CP-element group 405: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_update_completed_
      -- 
    ca_3100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => convTranspose_CP_39_elements(405)); -- 
    req_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => WPIPE_ConvTranspose_output_pipe_1348_inst_req_0); -- 
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_sample_completed_
      -- CP-element group 406: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_update_start_
      -- CP-element group 406: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Update/req
      -- 
    ack_3109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1348_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    req_3113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1348_inst_req_1); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_update_completed_
      -- CP-element group 407: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1348_Update/$exit
      -- 
    ack_3114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1348_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	403 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_sample_start_
      -- CP-element group 408: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Sample/req
      -- 
    req_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => WPIPE_ConvTranspose_output_pipe_1351_inst_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(403) & convTranspose_CP_39_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_sample_completed_
      -- CP-element group 409: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_update_start_
      -- CP-element group 409: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Sample/ack
      -- CP-element group 409: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Update/req
      -- 
    ack_3123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1351_inst_ack_0, ack => convTranspose_CP_39_elements(409)); -- 
    req_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1351_inst_req_1); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1351_Update/ack
      -- 
    ack_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1351_inst_ack_1, ack => convTranspose_CP_39_elements(410)); -- 
    -- CP-element group 411:  join  transition  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: 	401 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Sample/req
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_sample_start_
      -- 
    req_3136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => WPIPE_ConvTranspose_output_pipe_1354_inst_req_0); -- 
    convTranspose_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(410) & convTranspose_CP_39_elements(401);
      gj_convTranspose_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_update_start_
      -- CP-element group 412: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Update/req
      -- 
    ack_3137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1354_inst_ack_0, ack => convTranspose_CP_39_elements(412)); -- 
    req_3141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1354_inst_req_1); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1354_Update/ack
      -- 
    ack_3142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1354_inst_ack_1, ack => convTranspose_CP_39_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: 	399 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_sample_start_
      -- 
    req_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(414), ack => WPIPE_ConvTranspose_output_pipe_1357_inst_req_0); -- 
    convTranspose_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(413) & convTranspose_CP_39_elements(399);
      gj_convTranspose_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Update/req
      -- CP-element group 415: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Sample/ack
      -- CP-element group 415: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_update_start_
      -- CP-element group 415: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_sample_completed_
      -- 
    ack_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1357_inst_ack_0, ack => convTranspose_CP_39_elements(415)); -- 
    req_3155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1357_inst_req_1); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Update/ack
      -- CP-element group 416: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1357_update_completed_
      -- 
    ack_3156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1357_inst_ack_1, ack => convTranspose_CP_39_elements(416)); -- 
    -- CP-element group 417:  join  transition  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: 	397 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Sample/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_sample_start_
      -- 
    req_3164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => WPIPE_ConvTranspose_output_pipe_1360_inst_req_0); -- 
    convTranspose_cp_element_group_417: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_417"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(416) & convTranspose_CP_39_elements(397);
      gj_convTranspose_cp_element_group_417 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 418:  transition  input  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (6) 
      -- CP-element group 418: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Update/req
      -- CP-element group 418: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Sample/ack
      -- CP-element group 418: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_update_start_
      -- CP-element group 418: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_sample_completed_
      -- 
    ack_3165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1360_inst_ack_0, ack => convTranspose_CP_39_elements(418)); -- 
    req_3169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_ConvTranspose_output_pipe_1360_inst_req_1); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Update/ack
      -- CP-element group 419: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1360_update_completed_
      -- 
    ack_3170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1360_inst_ack_1, ack => convTranspose_CP_39_elements(419)); -- 
    -- CP-element group 420:  join  transition  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: 	395 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Sample/req
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_sample_start_
      -- 
    req_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(420), ack => WPIPE_ConvTranspose_output_pipe_1363_inst_req_0); -- 
    convTranspose_cp_element_group_420: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_420"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(419) & convTranspose_CP_39_elements(395);
      gj_convTranspose_cp_element_group_420 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 421:  transition  input  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (6) 
      -- CP-element group 421: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Update/req
      -- CP-element group 421: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Update/$entry
      -- CP-element group 421: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Sample/ack
      -- CP-element group 421: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_update_start_
      -- CP-element group 421: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_sample_completed_
      -- 
    ack_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1363_inst_ack_0, ack => convTranspose_CP_39_elements(421)); -- 
    req_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(421), ack => WPIPE_ConvTranspose_output_pipe_1363_inst_req_1); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Update/ack
      -- CP-element group 422: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1363_update_completed_
      -- 
    ack_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1363_inst_ack_1, ack => convTranspose_CP_39_elements(422)); -- 
    -- CP-element group 423:  join  transition  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: 	393 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Sample/req
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Sample/$entry
      -- CP-element group 423: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_sample_start_
      -- 
    req_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(423), ack => WPIPE_ConvTranspose_output_pipe_1366_inst_req_0); -- 
    convTranspose_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(422) & convTranspose_CP_39_elements(393);
      gj_convTranspose_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (6) 
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Update/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Sample/ack
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_sample_completed_
      -- 
    ack_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1366_inst_ack_0, ack => convTranspose_CP_39_elements(424)); -- 
    req_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => WPIPE_ConvTranspose_output_pipe_1366_inst_req_1); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_Update/ack
      -- CP-element group 425: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1366_update_completed_
      -- 
    ack_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1366_inst_ack_1, ack => convTranspose_CP_39_elements(425)); -- 
    -- CP-element group 426:  join  transition  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: 	391 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Sample/req
      -- 
    req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => WPIPE_ConvTranspose_output_pipe_1369_inst_req_0); -- 
    convTranspose_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(425) & convTranspose_CP_39_elements(391);
      gj_convTranspose_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (6) 
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_sample_completed_
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_update_start_
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Sample/ack
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Update/req
      -- CP-element group 427: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Update/$entry
      -- 
    ack_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1369_inst_ack_0, ack => convTranspose_CP_39_elements(427)); -- 
    req_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(427), ack => WPIPE_ConvTranspose_output_pipe_1369_inst_req_1); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Update/ack
      -- CP-element group 428: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/WPIPE_ConvTranspose_output_pipe_1369_Update/$exit
      -- 
    ack_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1369_inst_ack_1, ack => convTranspose_CP_39_elements(428)); -- 
    -- CP-element group 429:  branch  join  transition  place  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: 	384 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429: 	431 
    -- CP-element group 429:  members (10) 
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382__exit__
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383__entry__
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383_else_link/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383_if_link/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383_eval_test/branch_req
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383_eval_test/$exit
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383_eval_test/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/if_stmt_1383_dead_link/$entry
      -- CP-element group 429: 	 branch_block_stmt_33/R_exitcond1_1384_place
      -- CP-element group 429: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/$exit
      -- 
    branch_req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => if_stmt_1383_branch_req_0); -- 
    convTranspose_cp_element_group_429: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_429"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(428) & convTranspose_CP_39_elements(384);
      gj_convTranspose_cp_element_group_429 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(429), clk => clk, reset => reset); --
    end block;
    -- CP-element group 430:  merge  transition  place  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	459 
    -- CP-element group 430:  members (13) 
      -- CP-element group 430: 	 branch_block_stmt_33/merge_stmt_1389__exit__
      -- CP-element group 430: 	 branch_block_stmt_33/forx_xend438x_xloopexit_forx_xend438
      -- CP-element group 430: 	 branch_block_stmt_33/if_stmt_1383_if_link/if_choice_transition
      -- CP-element group 430: 	 branch_block_stmt_33/if_stmt_1383_if_link/$exit
      -- CP-element group 430: 	 branch_block_stmt_33/forx_xbody366_forx_xend438x_xloopexit
      -- CP-element group 430: 	 branch_block_stmt_33/forx_xbody366_forx_xend438x_xloopexit_PhiReq/$entry
      -- CP-element group 430: 	 branch_block_stmt_33/forx_xbody366_forx_xend438x_xloopexit_PhiReq/$exit
      -- CP-element group 430: 	 branch_block_stmt_33/merge_stmt_1389_PhiReqMerge
      -- CP-element group 430: 	 branch_block_stmt_33/merge_stmt_1389_PhiAck/$entry
      -- CP-element group 430: 	 branch_block_stmt_33/merge_stmt_1389_PhiAck/$exit
      -- CP-element group 430: 	 branch_block_stmt_33/merge_stmt_1389_PhiAck/dummy
      -- CP-element group 430: 	 branch_block_stmt_33/forx_xend438x_xloopexit_forx_xend438_PhiReq/$entry
      -- CP-element group 430: 	 branch_block_stmt_33/forx_xend438x_xloopexit_forx_xend438_PhiReq/$exit
      -- 
    if_choice_transition_3225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_1, ack => convTranspose_CP_39_elements(430)); -- 
    -- CP-element group 431:  fork  transition  place  input  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	429 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	454 
    -- CP-element group 431: 	455 
    -- CP-element group 431:  members (12) 
      -- CP-element group 431: 	 branch_block_stmt_33/if_stmt_1383_else_link/else_choice_transition
      -- CP-element group 431: 	 branch_block_stmt_33/if_stmt_1383_else_link/$exit
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Sample/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Sample/rr
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Update/$entry
      -- CP-element group 431: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_0, ack => convTranspose_CP_39_elements(431)); -- 
    rr_3504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(431), ack => type_cast_1261_inst_req_0); -- 
    cr_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(431), ack => type_cast_1261_inst_req_1); -- 
    -- CP-element group 432:  merge  branch  transition  place  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	120 
    -- CP-element group 432: 	165 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	121 
    -- CP-element group 432: 	122 
    -- CP-element group 432:  members (17) 
      -- CP-element group 432: 	 branch_block_stmt_33/merge_stmt_425__exit__
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_431__entry__
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_431__exit__
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432__entry__
      -- CP-element group 432: 	 branch_block_stmt_33/merge_stmt_425_PhiAck/dummy
      -- CP-element group 432: 	 branch_block_stmt_33/merge_stmt_425_PhiAck/$exit
      -- CP-element group 432: 	 branch_block_stmt_33/merge_stmt_425_PhiAck/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_431/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/assign_stmt_431/$exit
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432_dead_link/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432_eval_test/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432_eval_test/$exit
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432_eval_test/branch_req
      -- CP-element group 432: 	 branch_block_stmt_33/R_cmp194447_433_place
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432_if_link/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/if_stmt_432_else_link/$entry
      -- CP-element group 432: 	 branch_block_stmt_33/merge_stmt_425_PhiReqMerge
      -- 
    branch_req_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(432), ack => if_stmt_432_branch_req_0); -- 
    convTranspose_CP_39_elements(432) <= OrReduce(convTranspose_CP_39_elements(120) & convTranspose_CP_39_elements(165));
    -- CP-element group 433:  transition  output  delay-element  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	124 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	437 
    -- CP-element group 433:  members (5) 
      -- CP-element group 433: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_req
      -- CP-element group 433: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_474_konst_delay_trans
      -- CP-element group 433: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$exit
      -- CP-element group 433: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/phi_stmt_470/$exit
      -- CP-element group 433: 	 branch_block_stmt_33/bbx_xnph453_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_470_req_3277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_470_req_3277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(433), ack => phi_stmt_470_req_0); -- 
    -- Element group convTranspose_CP_39_elements(433) is a control-delay.
    cp_element_433_delay: control_delay_element  generic map(name => " 433_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(433), clk => clk, reset =>reset);
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	166 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	436 
    -- CP-element group 434:  members (2) 
      -- CP-element group 434: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Sample/ra
      -- 
    ra_3297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_476_inst_ack_0, ack => convTranspose_CP_39_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	166 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (2) 
      -- CP-element group 435: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/Update/ca
      -- 
    ca_3302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_476_inst_ack_1, ack => convTranspose_CP_39_elements(435)); -- 
    -- CP-element group 436:  join  transition  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	434 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (6) 
      -- CP-element group 436: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/SplitProtocol/$exit
      -- CP-element group 436: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_req
      -- CP-element group 436: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/type_cast_476/$exit
      -- CP-element group 436: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/phi_stmt_470_sources/$exit
      -- CP-element group 436: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_470/$exit
      -- CP-element group 436: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_470_req_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_470_req_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(436), ack => phi_stmt_470_req_1); -- 
    convTranspose_cp_element_group_436: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_436"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(434) & convTranspose_CP_39_elements(435);
      gj_convTranspose_cp_element_group_436 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(436), clk => clk, reset => reset); --
    end block;
    -- CP-element group 437:  merge  transition  place  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	433 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (2) 
      -- CP-element group 437: 	 branch_block_stmt_33/merge_stmt_469_PhiReqMerge
      -- CP-element group 437: 	 branch_block_stmt_33/merge_stmt_469_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(437) <= OrReduce(convTranspose_CP_39_elements(433) & convTranspose_CP_39_elements(436));
    -- CP-element group 438:  fork  transition  place  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	144 
    -- CP-element group 438: 	148 
    -- CP-element group 438: 	152 
    -- CP-element group 438: 	156 
    -- CP-element group 438: 	160 
    -- CP-element group 438: 	163 
    -- CP-element group 438: 	125 
    -- CP-element group 438: 	126 
    -- CP-element group 438: 	128 
    -- CP-element group 438: 	129 
    -- CP-element group 438: 	132 
    -- CP-element group 438: 	136 
    -- CP-element group 438: 	140 
    -- CP-element group 438:  members (56) 
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/merge_stmt_469__exit__
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632__entry__
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_575_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_557_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/word_0/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_539_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_593_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_611_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/ptr_deref_619_Update/word_access_complete/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resized_1
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scaled_1
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_computed_1
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/$exit
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/index_resize_req
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_resize_1/index_resize_ack
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/$exit
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/scale_rename_req
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_index_scale_1/scale_rename_ack
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_update_start
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Sample/req
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/array_obj_ref_482_final_index_sum_regn_Update/req
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/addr_of_483_complete/req
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_sample_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/RPIPE_ConvTranspose_input_pipe_486_Sample/rr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_490_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_503_Update/cr
      -- CP-element group 438: 	 branch_block_stmt_33/assign_stmt_484_to_assign_stmt_632/type_cast_521_update_start_
      -- CP-element group 438: 	 branch_block_stmt_33/merge_stmt_469_PhiAck/phi_stmt_470_ack
      -- CP-element group 438: 	 branch_block_stmt_33/merge_stmt_469_PhiAck/$exit
      -- 
    phi_stmt_470_ack_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_470_ack_0, ack => convTranspose_CP_39_elements(438)); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_575_inst_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_557_inst_req_1); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_521_inst_req_1); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_593_inst_req_1); -- 
    cr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => ptr_deref_619_store_0_req_1); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_539_inst_req_1); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_611_inst_req_1); -- 
    req_981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => array_obj_ref_482_index_offset_req_0); -- 
    req_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => array_obj_ref_482_index_offset_req_1); -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => addr_of_483_final_reg_req_1); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => RPIPE_ConvTranspose_input_pipe_486_inst_req_0); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_490_inst_req_1); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => type_cast_503_inst_req_1); -- 
    -- CP-element group 439:  transition  output  delay-element  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	168 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	443 
    -- CP-element group 439:  members (5) 
      -- CP-element group 439: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/$exit
      -- CP-element group 439: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/phi_stmt_677/$exit
      -- CP-element group 439: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_req
      -- CP-element group 439: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_681_konst_delay_trans
      -- CP-element group 439: 	 branch_block_stmt_33/bbx_xnph449_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$exit
      -- 
    phi_stmt_677_req_3331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_677_req_3331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(439), ack => phi_stmt_677_req_0); -- 
    -- Element group convTranspose_CP_39_elements(439) is a control-delay.
    cp_element_439_delay: control_delay_element  generic map(name => " 439_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(439), clk => clk, reset =>reset);
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	210 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	442 
    -- CP-element group 440:  members (2) 
      -- CP-element group 440: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/ra
      -- CP-element group 440: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Sample/$exit
      -- 
    ra_3351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_683_inst_ack_0, ack => convTranspose_CP_39_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	210 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (2) 
      -- CP-element group 441: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/ca
      -- CP-element group 441: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/Update/$exit
      -- 
    ca_3356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_683_inst_ack_1, ack => convTranspose_CP_39_elements(441)); -- 
    -- CP-element group 442:  join  transition  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	440 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (6) 
      -- CP-element group 442: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_req
      -- CP-element group 442: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/SplitProtocol/$exit
      -- CP-element group 442: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/type_cast_683/$exit
      -- CP-element group 442: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/phi_stmt_677_sources/$exit
      -- CP-element group 442: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_677/$exit
      -- CP-element group 442: 	 branch_block_stmt_33/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- 
    phi_stmt_677_req_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_677_req_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(442), ack => phi_stmt_677_req_1); -- 
    convTranspose_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(440) & convTranspose_CP_39_elements(441);
      gj_convTranspose_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  merge  transition  place  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	439 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (2) 
      -- CP-element group 443: 	 branch_block_stmt_33/merge_stmt_676_PhiReqMerge
      -- CP-element group 443: 	 branch_block_stmt_33/merge_stmt_676_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(443) <= OrReduce(convTranspose_CP_39_elements(439) & convTranspose_CP_39_elements(442));
    -- CP-element group 444:  fork  transition  place  input  output  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	184 
    -- CP-element group 444: 	188 
    -- CP-element group 444: 	192 
    -- CP-element group 444: 	196 
    -- CP-element group 444: 	200 
    -- CP-element group 444: 	204 
    -- CP-element group 444: 	180 
    -- CP-element group 444: 	207 
    -- CP-element group 444: 	169 
    -- CP-element group 444: 	170 
    -- CP-element group 444: 	172 
    -- CP-element group 444: 	173 
    -- CP-element group 444: 	176 
    -- CP-element group 444:  members (56) 
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_update_start
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_728_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/merge_stmt_676__exit__
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839__entry__
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_sample_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/scale_rename_ack
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/scale_rename_req
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/$exit
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scale_1/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_697_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_complete/req
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_710_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Update/req
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/index_resize_ack
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/index_resize_req
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/$exit
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resize_1/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_computed_1
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_scaled_1
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_index_resized_1
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/addr_of_690_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/req
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/rr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/array_obj_ref_689_final_index_sum_regn_Sample/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/RPIPE_ConvTranspose_input_pipe_693_Sample/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_746_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_764_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_782_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_800_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/type_cast_818_Update/cr
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_update_start_
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/$entry
      -- CP-element group 444: 	 branch_block_stmt_33/assign_stmt_691_to_assign_stmt_839/ptr_deref_826_Update/word_access_complete/word_0/cr
      -- CP-element group 444: 	 branch_block_stmt_33/merge_stmt_676_PhiAck/phi_stmt_677_ack
      -- CP-element group 444: 	 branch_block_stmt_33/merge_stmt_676_PhiAck/$exit
      -- 
    phi_stmt_677_ack_3362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_677_ack_0, ack => convTranspose_CP_39_elements(444)); -- 
    cr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_728_inst_req_1); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_697_inst_req_1); -- 
    req_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => addr_of_690_final_reg_req_1); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_710_inst_req_1); -- 
    req_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => array_obj_ref_689_index_offset_req_1); -- 
    req_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => array_obj_ref_689_index_offset_req_0); -- 
    rr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => RPIPE_ConvTranspose_input_pipe_693_inst_req_0); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_746_inst_req_1); -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_764_inst_req_1); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_782_inst_req_1); -- 
    cr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_800_inst_req_1); -- 
    cr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => type_cast_818_inst_req_1); -- 
    cr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => ptr_deref_826_store_0_req_1); -- 
    -- CP-element group 445:  merge  fork  transition  place  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	209 
    -- CP-element group 445: 	122 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	211 
    -- CP-element group 445: 	212 
    -- CP-element group 445: 	213 
    -- CP-element group 445: 	214 
    -- CP-element group 445: 	215 
    -- CP-element group 445: 	216 
    -- CP-element group 445:  members (25) 
      -- CP-element group 445: 	 branch_block_stmt_33/merge_stmt_848__exit__
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876__entry__
      -- CP-element group 445: 	 branch_block_stmt_33/merge_stmt_848_PhiReqMerge
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_update_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_851_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_update_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_855_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_update_start_
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_33/assign_stmt_852_to_assign_stmt_876/type_cast_859_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_33/merge_stmt_848_PhiAck/dummy
      -- CP-element group 445: 	 branch_block_stmt_33/merge_stmt_848_PhiAck/$exit
      -- CP-element group 445: 	 branch_block_stmt_33/merge_stmt_848_PhiAck/$entry
      -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => type_cast_851_inst_req_0); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => type_cast_851_inst_req_1); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => type_cast_855_inst_req_0); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => type_cast_855_inst_req_1); -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => type_cast_859_inst_req_0); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => type_cast_859_inst_req_1); -- 
    convTranspose_CP_39_elements(445) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 446:  transition  output  delay-element  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	221 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	450 
    -- CP-element group 446:  members (5) 
      -- CP-element group 446: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/phi_stmt_921/$exit
      -- CP-element group 446: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_927_konst_delay_trans
      -- CP-element group 446: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/$exit
      -- CP-element group 446: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$exit
      -- CP-element group 446: 	 branch_block_stmt_33/bbx_xnph445_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_req
      -- 
    phi_stmt_921_req_3408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_921_req_3408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(446), ack => phi_stmt_921_req_1); -- 
    -- Element group convTranspose_CP_39_elements(446) is a control-delay.
    cp_element_446_delay: control_delay_element  generic map(name => " 446_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(446), clk => clk, reset =>reset);
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	230 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	449 
    -- CP-element group 447:  members (2) 
      -- CP-element group 447: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Sample/ra
      -- 
    ra_3428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_0, ack => convTranspose_CP_39_elements(447)); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	230 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (2) 
      -- CP-element group 448: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/Update/ca
      -- 
    ca_3433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_1, ack => convTranspose_CP_39_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	447 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (6) 
      -- CP-element group 449: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_sources/type_cast_924/SplitProtocol/$exit
      -- CP-element group 449: 	 branch_block_stmt_33/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_921/phi_stmt_921_req
      -- 
    phi_stmt_921_req_3434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_921_req_3434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => phi_stmt_921_req_0); -- 
    convTranspose_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(447) & convTranspose_CP_39_elements(448);
      gj_convTranspose_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  merge  transition  place  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	446 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (2) 
      -- CP-element group 450: 	 branch_block_stmt_33/merge_stmt_920_PhiReqMerge
      -- CP-element group 450: 	 branch_block_stmt_33/merge_stmt_920_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(450) <= OrReduce(convTranspose_CP_39_elements(446) & convTranspose_CP_39_elements(449));
    -- CP-element group 451:  fork  transition  place  input  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	222 
    -- CP-element group 451: 	223 
    -- CP-element group 451: 	225 
    -- CP-element group 451: 	227 
    -- CP-element group 451:  members (29) 
      -- CP-element group 451: 	 branch_block_stmt_33/merge_stmt_920__exit__
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951__entry__
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_update_start_
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resized_1
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scaled_1
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_computed_1
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/$exit
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/index_resize_req
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_resize_1/index_resize_ack
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/$exit
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/scale_rename_req
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_index_scale_1/scale_rename_ack
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_update_start
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Sample/req
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/array_obj_ref_933_final_index_sum_regn_Update/req
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/addr_of_934_complete/req
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_update_start_
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/$entry
      -- CP-element group 451: 	 branch_block_stmt_33/assign_stmt_935_to_assign_stmt_951/ptr_deref_937_Update/word_access_complete/word_0/cr
      -- CP-element group 451: 	 branch_block_stmt_33/merge_stmt_920_PhiAck/$exit
      -- CP-element group 451: 	 branch_block_stmt_33/merge_stmt_920_PhiAck/phi_stmt_921_ack
      -- 
    phi_stmt_921_ack_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_921_ack_0, ack => convTranspose_CP_39_elements(451)); -- 
    req_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => array_obj_ref_933_index_offset_req_0); -- 
    req_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => array_obj_ref_933_index_offset_req_1); -- 
    req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => addr_of_934_final_reg_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => ptr_deref_937_store_0_req_1); -- 
    -- CP-element group 452:  merge  fork  transition  place  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	219 
    -- CP-element group 452: 	229 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	231 
    -- CP-element group 452: 	232 
    -- CP-element group 452: 	234 
    -- CP-element group 452: 	235 
    -- CP-element group 452: 	263 
    -- CP-element group 452: 	281 
    -- CP-element group 452: 	282 
    -- CP-element group 452: 	286 
    -- CP-element group 452: 	287 
    -- CP-element group 452: 	297 
    -- CP-element group 452: 	315 
    -- CP-element group 452: 	316 
    -- CP-element group 452: 	320 
    -- CP-element group 452: 	321 
    -- CP-element group 452: 	331 
    -- CP-element group 452: 	349 
    -- CP-element group 452: 	350 
    -- CP-element group 452: 	354 
    -- CP-element group 452: 	355 
    -- CP-element group 452: 	365 
    -- CP-element group 452: 	367 
    -- CP-element group 452: 	369 
    -- CP-element group 452: 	371 
    -- CP-element group 452:  members (76) 
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/merge_stmt_960__exit__
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193__entry__
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1056_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1043_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Sample/crr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/call_stmt_963_Update/ccr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_968_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1099_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1112_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1155_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_update_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/type_cast_1168_Update/cr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/call_stmt_963_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_33/merge_stmt_960_PhiReqMerge
      -- CP-element group 452: 	 branch_block_stmt_33/merge_stmt_960_PhiAck/$entry
      -- CP-element group 452: 	 branch_block_stmt_33/merge_stmt_960_PhiAck/$exit
      -- CP-element group 452: 	 branch_block_stmt_33/merge_stmt_960_PhiAck/dummy
      -- 
    rr_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1056_inst_req_0); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_Block1_start_1014_inst_req_0); -- 
    cr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1056_inst_req_1); -- 
    rr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1043_inst_req_0); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_Block2_start_1070_inst_req_0); -- 
    cr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1043_inst_req_1); -- 
    crr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => call_stmt_963_call_req_0); -- 
    ccr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => call_stmt_963_call_req_1); -- 
    cr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_968_inst_req_1); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_Block0_start_970_inst_req_0); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1099_inst_req_0); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1099_inst_req_1); -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1112_inst_req_0); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1112_inst_req_1); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_Block3_start_1126_inst_req_0); -- 
    rr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1155_inst_req_0); -- 
    cr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1155_inst_req_1); -- 
    rr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1168_inst_req_0); -- 
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => type_cast_1168_inst_req_1); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => RPIPE_Block0_done_1183_inst_req_0); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => RPIPE_Block1_done_1186_inst_req_0); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => RPIPE_Block2_done_1189_inst_req_0); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => RPIPE_Block3_done_1192_inst_req_0); -- 
    convTranspose_CP_39_elements(452) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 453:  transition  output  delay-element  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	383 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	457 
    -- CP-element group 453:  members (5) 
      -- CP-element group 453: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/$exit
      -- CP-element group 453: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/phi_stmt_1255/$exit
      -- CP-element group 453: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/$exit
      -- CP-element group 453: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1259_konst_delay_trans
      -- CP-element group 453: 	 branch_block_stmt_33/bbx_xnph_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_req
      -- 
    phi_stmt_1255_req_3485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1255_req_3485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(453), ack => phi_stmt_1255_req_0); -- 
    -- Element group convTranspose_CP_39_elements(453) is a control-delay.
    cp_element_453_delay: control_delay_element  generic map(name => " 453_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(383), ack => convTranspose_CP_39_elements(453), clk => clk, reset =>reset);
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	431 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (2) 
      -- CP-element group 454: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Sample/$exit
      -- CP-element group 454: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Sample/ra
      -- 
    ra_3505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_0, ack => convTranspose_CP_39_elements(454)); -- 
    -- CP-element group 455:  transition  input  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	431 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (2) 
      -- CP-element group 455: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Update/$exit
      -- CP-element group 455: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/Update/ca
      -- 
    ca_3510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_1, ack => convTranspose_CP_39_elements(455)); -- 
    -- CP-element group 456:  join  transition  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (6) 
      -- CP-element group 456: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_sources/type_cast_1261/SplitProtocol/$exit
      -- CP-element group 456: 	 branch_block_stmt_33/forx_xbody366_forx_xbody366_PhiReq/phi_stmt_1255/phi_stmt_1255_req
      -- 
    phi_stmt_1255_req_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1255_req_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => phi_stmt_1255_req_1); -- 
    convTranspose_cp_element_group_456: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_456"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(454) & convTranspose_CP_39_elements(455);
      gj_convTranspose_cp_element_group_456 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(456), clk => clk, reset => reset); --
    end block;
    -- CP-element group 457:  merge  transition  place  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	453 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (2) 
      -- CP-element group 457: 	 branch_block_stmt_33/merge_stmt_1254_PhiReqMerge
      -- CP-element group 457: 	 branch_block_stmt_33/merge_stmt_1254_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(457) <= OrReduce(convTranspose_CP_39_elements(453) & convTranspose_CP_39_elements(456));
    -- CP-element group 458:  fork  transition  place  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	403 
    -- CP-element group 458: 	405 
    -- CP-element group 458: 	384 
    -- CP-element group 458: 	385 
    -- CP-element group 458: 	387 
    -- CP-element group 458: 	389 
    -- CP-element group 458: 	391 
    -- CP-element group 458: 	393 
    -- CP-element group 458: 	395 
    -- CP-element group 458: 	397 
    -- CP-element group 458: 	399 
    -- CP-element group 458: 	401 
    -- CP-element group 458:  members (53) 
      -- CP-element group 458: 	 branch_block_stmt_33/merge_stmt_1254__exit__
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382__entry__
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1306_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/word_access_complete/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/word_access_complete/word_0/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_Update/word_access_complete/word_0/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1346_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1296_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1336_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1286_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1326_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1276_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/type_cast_1316_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_resized_1
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_scaled_1
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_computed_1
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_resize_1/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_resize_1/$exit
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_resize_1/index_resize_req
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_resize_1/index_resize_ack
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_scale_1/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_scale_1/$exit
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_scale_1/scale_rename_req
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_index_scale_1/scale_rename_ack
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_update_start
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Sample/req
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/array_obj_ref_1267_final_index_sum_regn_Update/req
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_complete/$entry
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/addr_of_1268_complete/req
      -- CP-element group 458: 	 branch_block_stmt_33/assign_stmt_1269_to_assign_stmt_1382/ptr_deref_1272_update_start_
      -- CP-element group 458: 	 branch_block_stmt_33/merge_stmt_1254_PhiAck/$exit
      -- CP-element group 458: 	 branch_block_stmt_33/merge_stmt_1254_PhiAck/phi_stmt_1255_ack
      -- 
    phi_stmt_1255_ack_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1255_ack_0, ack => convTranspose_CP_39_elements(458)); -- 
    cr_3043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1306_inst_req_1); -- 
    cr_3099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1346_inst_req_1); -- 
    cr_2982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => ptr_deref_1272_load_0_req_1); -- 
    cr_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1296_inst_req_1); -- 
    cr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1336_inst_req_1); -- 
    cr_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1286_inst_req_1); -- 
    cr_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1326_inst_req_1); -- 
    cr_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1276_inst_req_1); -- 
    cr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => type_cast_1316_inst_req_1); -- 
    req_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => array_obj_ref_1267_index_offset_req_0); -- 
    req_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => array_obj_ref_1267_index_offset_req_1); -- 
    req_2937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => addr_of_1268_final_reg_req_1); -- 
    -- CP-element group 459:  merge  transition  place  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	430 
    -- CP-element group 459: 	381 
    -- CP-element group 459: successors 
    -- CP-element group 459:  members (16) 
      -- CP-element group 459: 	 $exit
      -- CP-element group 459: 	 branch_block_stmt_33/$exit
      -- CP-element group 459: 	 branch_block_stmt_33/branch_block_stmt_33__exit__
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1391__exit__
      -- CP-element group 459: 	 branch_block_stmt_33/return__
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1393__exit__
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1391_PhiReqMerge
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1391_PhiAck/$entry
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1391_PhiAck/$exit
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1391_PhiAck/dummy
      -- CP-element group 459: 	 branch_block_stmt_33/return___PhiReq/$entry
      -- CP-element group 459: 	 branch_block_stmt_33/return___PhiReq/$exit
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1393_PhiReqMerge
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1393_PhiAck/$entry
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1393_PhiAck/$exit
      -- CP-element group 459: 	 branch_block_stmt_33/merge_stmt_1393_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(459) <= OrReduce(convTranspose_CP_39_elements(430) & convTranspose_CP_39_elements(381));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar463_932_resized : std_logic_vector(13 downto 0);
    signal R_indvar463_932_scaled : std_logic_vector(13 downto 0);
    signal R_indvar477_688_resized : std_logic_vector(10 downto 0);
    signal R_indvar477_688_scaled : std_logic_vector(10 downto 0);
    signal R_indvar493_481_resized : std_logic_vector(13 downto 0);
    signal R_indvar493_481_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1266_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1266_scaled : std_logic_vector(13 downto 0);
    signal add108_334 : std_logic_vector(15 downto 0);
    signal add117_359 : std_logic_vector(15 downto 0);
    signal add126_384 : std_logic_vector(15 downto 0);
    signal add12_83 : std_logic_vector(15 downto 0);
    signal add135_409 : std_logic_vector(15 downto 0);
    signal add150_509 : std_logic_vector(63 downto 0);
    signal add156_527 : std_logic_vector(63 downto 0);
    signal add162_545 : std_logic_vector(63 downto 0);
    signal add168_563 : std_logic_vector(63 downto 0);
    signal add174_581 : std_logic_vector(63 downto 0);
    signal add180_599 : std_logic_vector(63 downto 0);
    signal add186_617 : std_logic_vector(63 downto 0);
    signal add206_716 : std_logic_vector(63 downto 0);
    signal add212_734 : std_logic_vector(63 downto 0);
    signal add218_752 : std_logic_vector(63 downto 0);
    signal add21_108 : std_logic_vector(15 downto 0);
    signal add224_770 : std_logic_vector(63 downto 0);
    signal add230_788 : std_logic_vector(63 downto 0);
    signal add236_806 : std_logic_vector(63 downto 0);
    signal add242_824 : std_logic_vector(63 downto 0);
    signal add30_133 : std_logic_vector(15 downto 0);
    signal add39_158 : std_logic_vector(15 downto 0);
    signal add48_183 : std_logic_vector(15 downto 0);
    signal add57_208 : std_logic_vector(15 downto 0);
    signal add74_248 : std_logic_vector(31 downto 0);
    signal add79_253 : std_logic_vector(31 downto 0);
    signal add99_309 : std_logic_vector(15 downto 0);
    signal add_58 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1267_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1267_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1267_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1267_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1267_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1267_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_482_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_689_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_689_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_933_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_933_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_691 : std_logic_vector(31 downto 0);
    signal arrayidx269_935 : std_logic_vector(31 downto 0);
    signal arrayidx371_1269 : std_logic_vector(31 downto 0);
    signal arrayidx_484 : std_logic_vector(31 downto 0);
    signal call101_312 : std_logic_vector(7 downto 0);
    signal call106_325 : std_logic_vector(7 downto 0);
    signal call10_74 : std_logic_vector(7 downto 0);
    signal call110_337 : std_logic_vector(7 downto 0);
    signal call115_350 : std_logic_vector(7 downto 0);
    signal call119_362 : std_logic_vector(7 downto 0);
    signal call124_375 : std_logic_vector(7 downto 0);
    signal call128_387 : std_logic_vector(7 downto 0);
    signal call133_400 : std_logic_vector(7 downto 0);
    signal call143_487 : std_logic_vector(7 downto 0);
    signal call147_500 : std_logic_vector(7 downto 0);
    signal call14_86 : std_logic_vector(7 downto 0);
    signal call153_518 : std_logic_vector(7 downto 0);
    signal call159_536 : std_logic_vector(7 downto 0);
    signal call165_554 : std_logic_vector(7 downto 0);
    signal call171_572 : std_logic_vector(7 downto 0);
    signal call177_590 : std_logic_vector(7 downto 0);
    signal call183_608 : std_logic_vector(7 downto 0);
    signal call199_694 : std_logic_vector(7 downto 0);
    signal call19_99 : std_logic_vector(7 downto 0);
    signal call203_707 : std_logic_vector(7 downto 0);
    signal call209_725 : std_logic_vector(7 downto 0);
    signal call215_743 : std_logic_vector(7 downto 0);
    signal call221_761 : std_logic_vector(7 downto 0);
    signal call227_779 : std_logic_vector(7 downto 0);
    signal call233_797 : std_logic_vector(7 downto 0);
    signal call239_815 : std_logic_vector(7 downto 0);
    signal call23_111 : std_logic_vector(7 downto 0);
    signal call275_963 : std_logic_vector(63 downto 0);
    signal call28_124 : std_logic_vector(7 downto 0);
    signal call2_49 : std_logic_vector(7 downto 0);
    signal call32_136 : std_logic_vector(7 downto 0);
    signal call346_1184 : std_logic_vector(15 downto 0);
    signal call348_1187 : std_logic_vector(15 downto 0);
    signal call350_1190 : std_logic_vector(15 downto 0);
    signal call352_1193 : std_logic_vector(15 downto 0);
    signal call354_1196 : std_logic_vector(63 downto 0);
    signal call37_149 : std_logic_vector(7 downto 0);
    signal call41_161 : std_logic_vector(7 downto 0);
    signal call46_174 : std_logic_vector(7 downto 0);
    signal call50_186 : std_logic_vector(7 downto 0);
    signal call55_199 : std_logic_vector(7 downto 0);
    signal call5_61 : std_logic_vector(7 downto 0);
    signal call92_287 : std_logic_vector(7 downto 0);
    signal call97_300 : std_logic_vector(7 downto 0);
    signal call_36 : std_logic_vector(7 downto 0);
    signal cmp194447_431 : std_logic_vector(0 downto 0);
    signal cmp264443_876 : std_logic_vector(0 downto 0);
    signal cmp451_416 : std_logic_vector(0 downto 0);
    signal conv104_316 : std_logic_vector(15 downto 0);
    signal conv107_329 : std_logic_vector(15 downto 0);
    signal conv113_341 : std_logic_vector(15 downto 0);
    signal conv116_354 : std_logic_vector(15 downto 0);
    signal conv11_78 : std_logic_vector(15 downto 0);
    signal conv122_366 : std_logic_vector(15 downto 0);
    signal conv125_379 : std_logic_vector(15 downto 0);
    signal conv131_391 : std_logic_vector(15 downto 0);
    signal conv134_404 : std_logic_vector(15 downto 0);
    signal conv144_491 : std_logic_vector(63 downto 0);
    signal conv149_504 : std_logic_vector(63 downto 0);
    signal conv155_522 : std_logic_vector(63 downto 0);
    signal conv161_540 : std_logic_vector(63 downto 0);
    signal conv167_558 : std_logic_vector(63 downto 0);
    signal conv173_576 : std_logic_vector(63 downto 0);
    signal conv179_594 : std_logic_vector(63 downto 0);
    signal conv17_90 : std_logic_vector(15 downto 0);
    signal conv185_612 : std_logic_vector(63 downto 0);
    signal conv1_40 : std_logic_vector(15 downto 0);
    signal conv200_698 : std_logic_vector(63 downto 0);
    signal conv205_711 : std_logic_vector(63 downto 0);
    signal conv20_103 : std_logic_vector(15 downto 0);
    signal conv211_729 : std_logic_vector(63 downto 0);
    signal conv217_747 : std_logic_vector(63 downto 0);
    signal conv223_765 : std_logic_vector(63 downto 0);
    signal conv229_783 : std_logic_vector(63 downto 0);
    signal conv235_801 : std_logic_vector(63 downto 0);
    signal conv241_819 : std_logic_vector(63 downto 0);
    signal conv253_852 : std_logic_vector(31 downto 0);
    signal conv255_856 : std_logic_vector(31 downto 0);
    signal conv258_860 : std_logic_vector(31 downto 0);
    signal conv26_115 : std_logic_vector(15 downto 0);
    signal conv276_969 : std_logic_vector(63 downto 0);
    signal conv29_128 : std_logic_vector(15 downto 0);
    signal conv304_1044 : std_logic_vector(15 downto 0);
    signal conv307_1057 : std_logic_vector(15 downto 0);
    signal conv321_1100 : std_logic_vector(15 downto 0);
    signal conv324_1113 : std_logic_vector(15 downto 0);
    signal conv338_1156 : std_logic_vector(15 downto 0);
    signal conv341_1169 : std_logic_vector(15 downto 0);
    signal conv355_1201 : std_logic_vector(63 downto 0);
    signal conv35_140 : std_logic_vector(15 downto 0);
    signal conv375_1277 : std_logic_vector(7 downto 0);
    signal conv381_1287 : std_logic_vector(7 downto 0);
    signal conv387_1297 : std_logic_vector(7 downto 0);
    signal conv38_153 : std_logic_vector(15 downto 0);
    signal conv393_1307 : std_logic_vector(7 downto 0);
    signal conv399_1317 : std_logic_vector(7 downto 0);
    signal conv3_53 : std_logic_vector(15 downto 0);
    signal conv405_1327 : std_logic_vector(7 downto 0);
    signal conv411_1337 : std_logic_vector(7 downto 0);
    signal conv417_1347 : std_logic_vector(7 downto 0);
    signal conv44_165 : std_logic_vector(15 downto 0);
    signal conv47_178 : std_logic_vector(15 downto 0);
    signal conv53_190 : std_logic_vector(15 downto 0);
    signal conv56_203 : std_logic_vector(15 downto 0);
    signal conv61_212 : std_logic_vector(31 downto 0);
    signal conv63_216 : std_logic_vector(31 downto 0);
    signal conv65_220 : std_logic_vector(31 downto 0);
    signal conv82_257 : std_logic_vector(31 downto 0);
    signal conv84_261 : std_logic_vector(31 downto 0);
    signal conv87_265 : std_logic_vector(31 downto 0);
    signal conv8_65 : std_logic_vector(15 downto 0);
    signal conv90_269 : std_logic_vector(31 downto 0);
    signal conv95_291 : std_logic_vector(15 downto 0);
    signal conv98_304 : std_logic_vector(15 downto 0);
    signal exitcond1_1382 : std_logic_vector(0 downto 0);
    signal exitcond2_839 : std_logic_vector(0 downto 0);
    signal exitcond3_632 : std_logic_vector(0 downto 0);
    signal exitcond_951 : std_logic_vector(0 downto 0);
    signal iNsTr_14_242 : std_logic_vector(31 downto 0);
    signal iNsTr_180_1239 : std_logic_vector(63 downto 0);
    signal iNsTr_26_454 : std_logic_vector(63 downto 0);
    signal iNsTr_39_661 : std_logic_vector(63 downto 0);
    signal iNsTr_53_905 : std_logic_vector(63 downto 0);
    signal indvar463_921 : std_logic_vector(63 downto 0);
    signal indvar477_677 : std_logic_vector(63 downto 0);
    signal indvar493_470 : std_logic_vector(63 downto 0);
    signal indvar_1255 : std_logic_vector(63 downto 0);
    signal indvarx_xnext464_946 : std_logic_vector(63 downto 0);
    signal indvarx_xnext478_834 : std_logic_vector(63 downto 0);
    signal indvarx_xnext494_627 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1377 : std_logic_vector(63 downto 0);
    signal mul256_865 : std_logic_vector(31 downto 0);
    signal mul259_870 : std_logic_vector(31 downto 0);
    signal mul66_230 : std_logic_vector(31 downto 0);
    signal mul85_274 : std_logic_vector(31 downto 0);
    signal mul88_279 : std_logic_vector(31 downto 0);
    signal mul91_284 : std_logic_vector(31 downto 0);
    signal mul_225 : std_logic_vector(31 downto 0);
    signal ptr_deref_1272_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1272_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1272_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1272_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1272_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_619_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_619_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_619_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_619_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_619_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_619_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_826_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_826_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_826_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_826_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_826_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_826_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_937_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_937_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_937_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_937_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_937_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_937_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_322 : std_logic_vector(15 downto 0);
    signal shl114_347 : std_logic_vector(15 downto 0);
    signal shl123_372 : std_logic_vector(15 downto 0);
    signal shl132_397 : std_logic_vector(15 downto 0);
    signal shl146_497 : std_logic_vector(63 downto 0);
    signal shl152_515 : std_logic_vector(63 downto 0);
    signal shl158_533 : std_logic_vector(63 downto 0);
    signal shl164_551 : std_logic_vector(63 downto 0);
    signal shl170_569 : std_logic_vector(63 downto 0);
    signal shl176_587 : std_logic_vector(63 downto 0);
    signal shl182_605 : std_logic_vector(63 downto 0);
    signal shl18_96 : std_logic_vector(15 downto 0);
    signal shl202_704 : std_logic_vector(63 downto 0);
    signal shl208_722 : std_logic_vector(63 downto 0);
    signal shl214_740 : std_logic_vector(63 downto 0);
    signal shl220_758 : std_logic_vector(63 downto 0);
    signal shl226_776 : std_logic_vector(63 downto 0);
    signal shl232_794 : std_logic_vector(63 downto 0);
    signal shl238_812 : std_logic_vector(63 downto 0);
    signal shl27_121 : std_logic_vector(15 downto 0);
    signal shl36_146 : std_logic_vector(15 downto 0);
    signal shl45_171 : std_logic_vector(15 downto 0);
    signal shl54_196 : std_logic_vector(15 downto 0);
    signal shl96_297 : std_logic_vector(15 downto 0);
    signal shl9_71 : std_logic_vector(15 downto 0);
    signal shl_46 : std_logic_vector(15 downto 0);
    signal shr306_1053 : std_logic_vector(31 downto 0);
    signal shr323_1109 : std_logic_vector(31 downto 0);
    signal shr340_1165 : std_logic_vector(31 downto 0);
    signal shr378_1283 : std_logic_vector(63 downto 0);
    signal shr384_1293 : std_logic_vector(63 downto 0);
    signal shr390_1303 : std_logic_vector(63 downto 0);
    signal shr396_1313 : std_logic_vector(63 downto 0);
    signal shr402_1323 : std_logic_vector(63 downto 0);
    signal shr408_1333 : std_logic_vector(63 downto 0);
    signal shr414_1343 : std_logic_vector(63 downto 0);
    signal shr_236 : std_logic_vector(31 downto 0);
    signal sub_1206 : std_logic_vector(63 downto 0);
    signal tmp372_1273 : std_logic_vector(63 downto 0);
    signal tmp458_1223 : std_logic_vector(31 downto 0);
    signal tmp458x_xop_1235 : std_logic_vector(31 downto 0);
    signal tmp459_1229 : std_logic_vector(0 downto 0);
    signal tmp462_1252 : std_logic_vector(63 downto 0);
    signal tmp470_889 : std_logic_vector(31 downto 0);
    signal tmp470x_xop_901 : std_logic_vector(31 downto 0);
    signal tmp471_895 : std_logic_vector(0 downto 0);
    signal tmp475_918 : std_logic_vector(63 downto 0);
    signal tmp486_645 : std_logic_vector(31 downto 0);
    signal tmp486x_xop_657 : std_logic_vector(31 downto 0);
    signal tmp487_651 : std_logic_vector(0 downto 0);
    signal tmp491_674 : std_logic_vector(63 downto 0);
    signal tmp500x_xop_450 : std_logic_vector(31 downto 0);
    signal tmp501_444 : std_logic_vector(0 downto 0);
    signal tmp505_467 : std_logic_vector(63 downto 0);
    signal type_cast_1003_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1051_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1107_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1199_wire : std_logic_vector(63 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1221_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1250_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1259_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1261_wire : std_logic_vector(63 downto 0);
    signal type_cast_1281_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1291_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1301_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1321_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1331_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1341_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1375_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_169_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_234_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_240_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_295_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_345_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_370_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_395_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_413_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_442_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_44_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_465_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_476_wire : std_logic_vector(63 downto 0);
    signal type_cast_495_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_531_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_585_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_603_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_625_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_643_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_655_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_672_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_681_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_683_wire : std_logic_vector(63 downto 0);
    signal type_cast_69_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_702_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_792_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_810_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_832_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_887_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_899_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_909_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_916_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_924_wire : std_logic_vector(63 downto 0);
    signal type_cast_927_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_939_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_967_wire : std_logic_vector(63 downto 0);
    signal type_cast_999_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop507_911 : std_logic_vector(63 downto 0);
    signal xx_xop508_667 : std_logic_vector(63 downto 0);
    signal xx_xop509_460 : std_logic_vector(63 downto 0);
    signal xx_xop_1245 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1267_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1267_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1267_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1267_resized_base_address <= "00000000000000";
    array_obj_ref_482_constant_part_of_offset <= "00000000000000";
    array_obj_ref_482_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_482_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_482_resized_base_address <= "00000000000000";
    array_obj_ref_689_constant_part_of_offset <= "00000100010";
    array_obj_ref_689_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_689_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_689_resized_base_address <= "00000000000";
    array_obj_ref_933_constant_part_of_offset <= "00000000000000";
    array_obj_ref_933_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_933_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_933_resized_base_address <= "00000000000000";
    ptr_deref_1272_word_offset_0 <= "00000000000000";
    ptr_deref_619_word_offset_0 <= "00000000000000";
    ptr_deref_826_word_offset_0 <= "00000000000";
    ptr_deref_937_word_offset_0 <= "00000000000000";
    type_cast_1003_wire_constant <= "0000000000000000";
    type_cast_1051_wire_constant <= "00000000000000000000000000010010";
    type_cast_1107_wire_constant <= "00000000000000000000000000010001";
    type_cast_1163_wire_constant <= "00000000000000000000000000010000";
    type_cast_119_wire_constant <= "0000000000001000";
    type_cast_1221_wire_constant <= "00000000000000000000000000000010";
    type_cast_1227_wire_constant <= "00000000000000000000000000000001";
    type_cast_1233_wire_constant <= "11111111111111111111111111111111";
    type_cast_1243_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1250_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1259_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1281_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1291_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1301_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1321_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1331_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1341_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1375_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_144_wire_constant <= "0000000000001000";
    type_cast_169_wire_constant <= "0000000000001000";
    type_cast_194_wire_constant <= "0000000000001000";
    type_cast_234_wire_constant <= "00000000000000000000000000000010";
    type_cast_240_wire_constant <= "00000000000000000000000000000001";
    type_cast_246_wire_constant <= "01111111111111111111111111111110";
    type_cast_295_wire_constant <= "0000000000001000";
    type_cast_320_wire_constant <= "0000000000001000";
    type_cast_345_wire_constant <= "0000000000001000";
    type_cast_370_wire_constant <= "0000000000001000";
    type_cast_395_wire_constant <= "0000000000001000";
    type_cast_413_wire_constant <= "00000000000000000000000000000011";
    type_cast_429_wire_constant <= "00000000000000000000000000000011";
    type_cast_442_wire_constant <= "00000000000000000000000000000001";
    type_cast_448_wire_constant <= "11111111111111111111111111111111";
    type_cast_44_wire_constant <= "0000000000001000";
    type_cast_458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_465_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_474_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_495_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_531_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_603_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_625_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_643_wire_constant <= "00000000000000000000000000000010";
    type_cast_649_wire_constant <= "00000000000000000000000000000001";
    type_cast_655_wire_constant <= "11111111111111111111111111111111";
    type_cast_665_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_672_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_681_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_69_wire_constant <= "0000000000001000";
    type_cast_702_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_720_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_738_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_792_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_810_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_832_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_874_wire_constant <= "00000000000000000000000000000011";
    type_cast_887_wire_constant <= "00000000000000000000000000000010";
    type_cast_893_wire_constant <= "00000000000000000000000000000001";
    type_cast_899_wire_constant <= "11111111111111111111111111111111";
    type_cast_909_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_916_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_927_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_939_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_944_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_94_wire_constant <= "0000000000001000";
    type_cast_999_wire_constant <= "0000000000000000";
    phi_stmt_1255: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1259_wire_constant & type_cast_1261_wire;
      req <= phi_stmt_1255_req_0 & phi_stmt_1255_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1255",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1255_ack_0,
          idata => idata,
          odata => indvar_1255,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1255
    phi_stmt_470: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_474_wire_constant & type_cast_476_wire;
      req <= phi_stmt_470_req_0 & phi_stmt_470_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_470",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_470_ack_0,
          idata => idata,
          odata => indvar493_470,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_470
    phi_stmt_677: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_681_wire_constant & type_cast_683_wire;
      req <= phi_stmt_677_req_0 & phi_stmt_677_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_677",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_677_ack_0,
          idata => idata,
          odata => indvar477_677,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_677
    phi_stmt_921: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_924_wire & type_cast_927_wire_constant;
      req <= phi_stmt_921_req_0 & phi_stmt_921_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_921",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_921_ack_0,
          idata => idata,
          odata => indvar463_921,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_921
    -- flow-through select operator MUX_1251_inst
    tmp462_1252 <= xx_xop_1245 when (tmp459_1229(0) /=  '0') else type_cast_1250_wire_constant;
    -- flow-through select operator MUX_466_inst
    tmp505_467 <= xx_xop509_460 when (tmp501_444(0) /=  '0') else type_cast_465_wire_constant;
    -- flow-through select operator MUX_673_inst
    tmp491_674 <= xx_xop508_667 when (tmp487_651(0) /=  '0') else type_cast_672_wire_constant;
    -- flow-through select operator MUX_917_inst
    tmp475_918 <= xx_xop507_911 when (tmp471_895(0) /=  '0') else type_cast_916_wire_constant;
    addr_of_1268_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1268_final_reg_req_0;
      addr_of_1268_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1268_final_reg_req_1;
      addr_of_1268_final_reg_ack_1<= rack(0);
      addr_of_1268_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1268_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1267_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx371_1269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_483_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_483_final_reg_req_0;
      addr_of_483_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_483_final_reg_req_1;
      addr_of_483_final_reg_ack_1<= rack(0);
      addr_of_483_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_483_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_482_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_690_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_690_final_reg_req_0;
      addr_of_690_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_690_final_reg_req_1;
      addr_of_690_final_reg_ack_1<= rack(0);
      addr_of_690_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_690_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_689_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_691,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_934_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_934_final_reg_req_0;
      addr_of_934_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_934_final_reg_req_1;
      addr_of_934_final_reg_ack_1<= rack(0);
      addr_of_934_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_934_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_933_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_102_inst_req_0;
      type_cast_102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_102_inst_req_1;
      type_cast_102_inst_ack_1<= rack(0);
      type_cast_102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1043_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1043_inst_req_0;
      type_cast_1043_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1043_inst_req_1;
      type_cast_1043_inst_ack_1<= rack(0);
      type_cast_1043_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1043_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_1044,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1056_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1056_inst_req_0;
      type_cast_1056_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1056_inst_req_1;
      type_cast_1056_inst_ack_1<= rack(0);
      type_cast_1056_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1056_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr306_1053,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1099_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1099_inst_req_0;
      type_cast_1099_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1099_inst_req_1;
      type_cast_1099_inst_ack_1<= rack(0);
      type_cast_1099_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1099_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv321_1100,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1112_inst_req_0;
      type_cast_1112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1112_inst_req_1;
      type_cast_1112_inst_ack_1<= rack(0);
      type_cast_1112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr323_1109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_114_inst_req_0;
      type_cast_114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_114_inst_req_1;
      type_cast_114_inst_ack_1<= rack(0);
      type_cast_114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1155_inst_req_0;
      type_cast_1155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1155_inst_req_1;
      type_cast_1155_inst_ack_1<= rack(0);
      type_cast_1155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv338_1156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1168_inst_req_0;
      type_cast_1168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1168_inst_req_1;
      type_cast_1168_inst_ack_1<= rack(0);
      type_cast_1168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr340_1165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1200_inst_req_0;
      type_cast_1200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1200_inst_req_1;
      type_cast_1200_inst_ack_1<= rack(0);
      type_cast_1200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1199_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp458x_xop_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_180_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1261_inst_req_0;
      type_cast_1261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1261_inst_req_1;
      type_cast_1261_inst_ack_1<= rack(0);
      type_cast_1261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1261_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1276_inst_req_0;
      type_cast_1276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1276_inst_req_1;
      type_cast_1276_inst_ack_1<= rack(0);
      type_cast_1276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp372_1273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv375_1277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_127_inst_req_0;
      type_cast_127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_127_inst_req_1;
      type_cast_127_inst_ack_1<= rack(0);
      type_cast_127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1286_inst_req_0;
      type_cast_1286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1286_inst_req_1;
      type_cast_1286_inst_ack_1<= rack(0);
      type_cast_1286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr378_1283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv381_1287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1296_inst_req_0;
      type_cast_1296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1296_inst_req_1;
      type_cast_1296_inst_ack_1<= rack(0);
      type_cast_1296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1296_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr384_1293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv387_1297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1306_inst_req_0;
      type_cast_1306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1306_inst_req_1;
      type_cast_1306_inst_ack_1<= rack(0);
      type_cast_1306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr390_1303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv393_1307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1316_inst_req_0;
      type_cast_1316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1316_inst_req_1;
      type_cast_1316_inst_ack_1<= rack(0);
      type_cast_1316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr396_1313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv399_1317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1326_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1326_inst_req_0;
      type_cast_1326_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1326_inst_req_1;
      type_cast_1326_inst_ack_1<= rack(0);
      type_cast_1326_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1326_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr402_1323,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv405_1327,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1336_inst_req_0;
      type_cast_1336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1336_inst_req_1;
      type_cast_1336_inst_ack_1<= rack(0);
      type_cast_1336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr408_1333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr414_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv417_1347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_152_inst_req_0;
      type_cast_152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_152_inst_req_1;
      type_cast_152_inst_ack_1<= rack(0);
      type_cast_152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_177_inst_req_0;
      type_cast_177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_177_inst_req_1;
      type_cast_177_inst_ack_1<= rack(0);
      type_cast_177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_189_inst_req_0;
      type_cast_189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_189_inst_req_1;
      type_cast_189_inst_ack_1<= rack(0);
      type_cast_189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_202_inst_req_0;
      type_cast_202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_202_inst_req_1;
      type_cast_202_inst_ack_1<= rack(0);
      type_cast_202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_58,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_215_inst_req_0;
      type_cast_215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_215_inst_req_1;
      type_cast_215_inst_ack_1<= rack(0);
      type_cast_215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_83,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_256_inst_req_0;
      type_cast_256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_256_inst_req_1;
      type_cast_256_inst_ack_1<= rack(0);
      type_cast_256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_260_inst_req_0;
      type_cast_260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_260_inst_req_1;
      type_cast_260_inst_ack_1<= rack(0);
      type_cast_260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_264_inst_req_0;
      type_cast_264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_264_inst_req_1;
      type_cast_264_inst_ack_1<= rack(0);
      type_cast_264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_265,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_268_inst_req_0;
      type_cast_268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_268_inst_req_1;
      type_cast_268_inst_ack_1<= rack(0);
      type_cast_268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_290_inst_req_0;
      type_cast_290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_290_inst_req_1;
      type_cast_290_inst_ack_1<= rack(0);
      type_cast_290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_303_inst_req_0;
      type_cast_303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_303_inst_req_1;
      type_cast_303_inst_ack_1<= rack(0);
      type_cast_303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_315_inst_req_0;
      type_cast_315_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_315_inst_req_1;
      type_cast_315_inst_ack_1<= rack(0);
      type_cast_315_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_316,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_328_inst_req_0;
      type_cast_328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_328_inst_req_1;
      type_cast_328_inst_ack_1<= rack(0);
      type_cast_328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_340_inst_req_0;
      type_cast_340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_340_inst_req_1;
      type_cast_340_inst_ack_1<= rack(0);
      type_cast_340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_353_inst_req_0;
      type_cast_353_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_353_inst_req_1;
      type_cast_353_inst_ack_1<= rack(0);
      type_cast_353_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_353_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_365_inst_req_0;
      type_cast_365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_365_inst_req_1;
      type_cast_365_inst_ack_1<= rack(0);
      type_cast_365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_378_inst_req_0;
      type_cast_378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_378_inst_req_1;
      type_cast_378_inst_ack_1<= rack(0);
      type_cast_378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_390_inst_req_0;
      type_cast_390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_390_inst_req_1;
      type_cast_390_inst_ack_1<= rack(0);
      type_cast_390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_39_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_39_inst_req_0;
      type_cast_39_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_39_inst_req_1;
      type_cast_39_inst_ack_1<= rack(0);
      type_cast_39_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_39_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_40,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_403_inst_req_0;
      type_cast_403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_403_inst_req_1;
      type_cast_403_inst_ack_1<= rack(0);
      type_cast_403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_400,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_404,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_453_inst_req_0;
      type_cast_453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_453_inst_req_1;
      type_cast_453_inst_ack_1<= rack(0);
      type_cast_453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_453_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp500x_xop_450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_476_inst_req_0;
      type_cast_476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_476_inst_req_1;
      type_cast_476_inst_ack_1<= rack(0);
      type_cast_476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext494_627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_476_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_490_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_490_inst_req_0;
      type_cast_490_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_490_inst_req_1;
      type_cast_490_inst_ack_1<= rack(0);
      type_cast_490_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_490_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_491,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_503_inst_req_0;
      type_cast_503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_503_inst_req_1;
      type_cast_503_inst_ack_1<= rack(0);
      type_cast_503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_521_inst_req_0;
      type_cast_521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_521_inst_req_1;
      type_cast_521_inst_ack_1<= rack(0);
      type_cast_521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_52_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_52_inst_req_0;
      type_cast_52_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_52_inst_req_1;
      type_cast_52_inst_ack_1<= rack(0);
      type_cast_52_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_52_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_539_inst_req_0;
      type_cast_539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_539_inst_req_1;
      type_cast_539_inst_ack_1<= rack(0);
      type_cast_539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_557_inst_req_0;
      type_cast_557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_557_inst_req_1;
      type_cast_557_inst_ack_1<= rack(0);
      type_cast_557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_575_inst_req_0;
      type_cast_575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_575_inst_req_1;
      type_cast_575_inst_ack_1<= rack(0);
      type_cast_575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_576,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_611_inst_req_0;
      type_cast_611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_611_inst_req_1;
      type_cast_611_inst_ack_1<= rack(0);
      type_cast_611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_61,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_65,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_660_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_660_inst_req_0;
      type_cast_660_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_660_inst_req_1;
      type_cast_660_inst_ack_1<= rack(0);
      type_cast_660_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_660_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp486x_xop_657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_683_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_683_inst_req_0;
      type_cast_683_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_683_inst_req_1;
      type_cast_683_inst_ack_1<= rack(0);
      type_cast_683_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_683_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext478_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_683_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_697_inst_req_0;
      type_cast_697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_697_inst_req_1;
      type_cast_697_inst_ack_1<= rack(0);
      type_cast_697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_710_inst_req_0;
      type_cast_710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_710_inst_req_1;
      type_cast_710_inst_ack_1<= rack(0);
      type_cast_710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_707,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_728_inst_req_0;
      type_cast_728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_728_inst_req_1;
      type_cast_728_inst_ack_1<= rack(0);
      type_cast_728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_746_inst_req_0;
      type_cast_746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_746_inst_req_1;
      type_cast_746_inst_ack_1<= rack(0);
      type_cast_746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_747,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_764_inst_req_0;
      type_cast_764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_764_inst_req_1;
      type_cast_764_inst_ack_1<= rack(0);
      type_cast_764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_77_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_77_inst_req_0;
      type_cast_77_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_77_inst_req_1;
      type_cast_77_inst_ack_1<= rack(0);
      type_cast_77_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_77_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_74,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_78,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_782_inst_req_0;
      type_cast_782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_782_inst_req_1;
      type_cast_782_inst_ack_1<= rack(0);
      type_cast_782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_800_inst_req_0;
      type_cast_800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_800_inst_req_1;
      type_cast_800_inst_ack_1<= rack(0);
      type_cast_800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_818_inst_req_0;
      type_cast_818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_818_inst_req_1;
      type_cast_818_inst_ack_1<= rack(0);
      type_cast_818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_818_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_819,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_359,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_855_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_855_inst_req_0;
      type_cast_855_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_855_inst_req_1;
      type_cast_855_inst_ack_1<= rack(0);
      type_cast_855_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_855_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_859_inst_req_0;
      type_cast_859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_859_inst_req_1;
      type_cast_859_inst_ack_1<= rack(0);
      type_cast_859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_89_inst_req_0;
      type_cast_89_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_89_inst_req_1;
      type_cast_89_inst_ack_1<= rack(0);
      type_cast_89_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_89_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_90,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_904_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_904_inst_req_0;
      type_cast_904_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_904_inst_req_1;
      type_cast_904_inst_ack_1<= rack(0);
      type_cast_904_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_904_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp470x_xop_901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_905,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_924_inst_req_0;
      type_cast_924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_924_inst_req_1;
      type_cast_924_inst_ack_1<= rack(0);
      type_cast_924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext464_946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_924_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_968_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_968_inst_req_0;
      type_cast_968_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_968_inst_req_1;
      type_cast_968_inst_ack_1<= rack(0);
      type_cast_968_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_968_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_967_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_969,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1267_index_1_rename
    process(R_indvar_1266_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1266_resized;
      ov(13 downto 0) := iv;
      R_indvar_1266_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1267_index_1_resize
    process(indvar_1255) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1255;
      ov := iv(13 downto 0);
      R_indvar_1266_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1267_root_address_inst
    process(array_obj_ref_1267_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1267_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1267_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_482_index_1_rename
    process(R_indvar493_481_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar493_481_resized;
      ov(13 downto 0) := iv;
      R_indvar493_481_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_482_index_1_resize
    process(indvar493_470) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar493_470;
      ov := iv(13 downto 0);
      R_indvar493_481_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_482_root_address_inst
    process(array_obj_ref_482_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_482_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_482_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_689_index_1_rename
    process(R_indvar477_688_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar477_688_resized;
      ov(10 downto 0) := iv;
      R_indvar477_688_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_689_index_1_resize
    process(indvar477_677) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar477_677;
      ov := iv(10 downto 0);
      R_indvar477_688_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_689_root_address_inst
    process(array_obj_ref_689_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_689_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_689_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_933_index_1_rename
    process(R_indvar463_932_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar463_932_resized;
      ov(13 downto 0) := iv;
      R_indvar463_932_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_933_index_1_resize
    process(indvar463_921) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar463_921;
      ov := iv(13 downto 0);
      R_indvar463_932_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_933_root_address_inst
    process(array_obj_ref_933_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_933_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_933_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1272_addr_0
    process(ptr_deref_1272_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1272_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1272_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1272_base_resize
    process(arrayidx371_1269) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx371_1269;
      ov := iv(13 downto 0);
      ptr_deref_1272_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1272_gather_scatter
    process(ptr_deref_1272_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1272_data_0;
      ov(63 downto 0) := iv;
      tmp372_1273 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1272_root_address_inst
    process(ptr_deref_1272_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1272_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1272_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_addr_0
    process(ptr_deref_619_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_619_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_619_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_base_resize
    process(arrayidx_484) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_484;
      ov := iv(13 downto 0);
      ptr_deref_619_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_gather_scatter
    process(add186_617) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_617;
      ov(63 downto 0) := iv;
      ptr_deref_619_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_619_root_address_inst
    process(ptr_deref_619_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_619_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_619_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_addr_0
    process(ptr_deref_826_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_826_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_826_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_base_resize
    process(arrayidx246_691) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_691;
      ov := iv(10 downto 0);
      ptr_deref_826_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_gather_scatter
    process(add242_824) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_824;
      ov(63 downto 0) := iv;
      ptr_deref_826_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_826_root_address_inst
    process(ptr_deref_826_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_826_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_826_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_addr_0
    process(ptr_deref_937_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_937_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_937_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_base_resize
    process(arrayidx269_935) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_935;
      ov := iv(13 downto 0);
      ptr_deref_937_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_gather_scatter
    process(type_cast_939_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_939_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_937_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_937_root_address_inst
    process(ptr_deref_937_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_937_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_937_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1211_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264443_876;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1211_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1211_branch_req_0,
          ack0 => if_stmt_1211_branch_ack_0,
          ack1 => if_stmt_1211_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1383_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1382;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1383_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1383_branch_req_0,
          ack0 => if_stmt_1383_branch_ack_0,
          ack1 => if_stmt_1383_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_417_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp451_416;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_417_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_417_branch_req_0,
          ack0 => if_stmt_417_branch_ack_0,
          ack1 => if_stmt_417_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_432_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194447_431;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_432_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_432_branch_req_0,
          ack0 => if_stmt_432_branch_ack_0,
          ack1 => if_stmt_432_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_633_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_632;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_633_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_633_branch_req_0,
          ack0 => if_stmt_633_branch_ack_0,
          ack1 => if_stmt_633_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_840_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_839;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_840_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_840_branch_req_0,
          ack0 => if_stmt_840_branch_ack_0,
          ack1 => if_stmt_840_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_877_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264443_876;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_877_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_877_branch_req_0,
          ack0 => if_stmt_877_branch_ack_0,
          ack1 => if_stmt_877_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_952_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_951;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_952_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_952_branch_req_0,
          ack0 => if_stmt_952_branch_ack_0,
          ack1 => if_stmt_952_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1234_inst
    process(tmp458_1223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp458_1223, type_cast_1233_wire_constant, tmp_var);
      tmp458x_xop_1235 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_252_inst
    process(add74_248, shr_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_248, shr_236, tmp_var);
      add79_253 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_449_inst
    process(shr_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_236, type_cast_448_wire_constant, tmp_var);
      tmp500x_xop_450 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_656_inst
    process(tmp486_645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp486_645, type_cast_655_wire_constant, tmp_var);
      tmp486x_xop_657 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_900_inst
    process(tmp470_889) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp470_889, type_cast_899_wire_constant, tmp_var);
      tmp470x_xop_901 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1244_inst
    process(iNsTr_180_1239) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_180_1239, type_cast_1243_wire_constant, tmp_var);
      xx_xop_1245 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1376_inst
    process(indvar_1255) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1255, type_cast_1375_wire_constant, tmp_var);
      indvarx_xnext_1377 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_459_inst
    process(iNsTr_26_454) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_454, type_cast_458_wire_constant, tmp_var);
      xx_xop509_460 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_626_inst
    process(indvar493_470) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar493_470, type_cast_625_wire_constant, tmp_var);
      indvarx_xnext494_627 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_666_inst
    process(iNsTr_39_661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_661, type_cast_665_wire_constant, tmp_var);
      xx_xop508_667 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_833_inst
    process(indvar477_677) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar477_677, type_cast_832_wire_constant, tmp_var);
      indvarx_xnext478_834 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_910_inst
    process(iNsTr_53_905) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_905, type_cast_909_wire_constant, tmp_var);
      xx_xop507_911 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_945_inst
    process(indvar463_921) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar463_921, type_cast_944_wire_constant, tmp_var);
      indvarx_xnext464_946 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_247_inst
    process(iNsTr_14_242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_242, type_cast_246_wire_constant, tmp_var);
      add74_248 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1381_inst
    process(indvarx_xnext_1377, tmp462_1252) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1377, tmp462_1252, tmp_var);
      exitcond1_1382 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_631_inst
    process(indvarx_xnext494_627, tmp505_467) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext494_627, tmp505_467, tmp_var);
      exitcond3_632 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_838_inst
    process(indvarx_xnext478_834, tmp491_674) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext478_834, tmp491_674, tmp_var);
      exitcond2_839 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_950_inst
    process(indvarx_xnext464_946, tmp475_918) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext464_946, tmp475_918, tmp_var);
      exitcond_951 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1052_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_1051_wire_constant, tmp_var);
      shr306_1053 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1108_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_1107_wire_constant, tmp_var);
      shr323_1109 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1164_inst
    process(add79_253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_253, type_cast_1163_wire_constant, tmp_var);
      shr340_1165 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1222_inst
    process(mul259_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_870, type_cast_1221_wire_constant, tmp_var);
      tmp458_1223 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_235_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_234_wire_constant, tmp_var);
      shr_236 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_241_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_240_wire_constant, tmp_var);
      iNsTr_14_242 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_644_inst
    process(mul91_284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_284, type_cast_643_wire_constant, tmp_var);
      tmp486_645 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_888_inst
    process(mul259_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_870, type_cast_887_wire_constant, tmp_var);
      tmp470_889 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1282_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1281_wire_constant, tmp_var);
      shr378_1283 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1292_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1291_wire_constant, tmp_var);
      shr384_1293 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1302_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1301_wire_constant, tmp_var);
      shr390_1303 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1312_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1311_wire_constant, tmp_var);
      shr396_1313 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1322_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1321_wire_constant, tmp_var);
      shr402_1323 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1332_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1331_wire_constant, tmp_var);
      shr408_1333 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1342_inst
    process(tmp372_1273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp372_1273, type_cast_1341_wire_constant, tmp_var);
      shr414_1343 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_224_inst
    process(conv63_216, conv61_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_216, conv61_212, tmp_var);
      mul_225 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(mul_225, conv65_220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_225, conv65_220, tmp_var);
      mul66_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_273_inst
    process(conv84_261, conv82_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_261, conv82_257, tmp_var);
      mul85_274 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_278_inst
    process(mul85_274, conv87_265) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_274, conv87_265, tmp_var);
      mul88_279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_283_inst
    process(mul88_279, conv90_269) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_279, conv90_269, tmp_var);
      mul91_284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_864_inst
    process(conv255_856, conv253_852) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_856, conv253_852, tmp_var);
      mul256_865 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_869_inst
    process(mul256_865, conv258_860) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_865, conv258_860, tmp_var);
      mul259_870 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_107_inst
    process(shl18_96, conv20_103) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_96, conv20_103, tmp_var);
      add21_108 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_132_inst
    process(shl27_121, conv29_128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_121, conv29_128, tmp_var);
      add30_133 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_157_inst
    process(shl36_146, conv38_153) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_146, conv38_153, tmp_var);
      add39_158 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_182_inst
    process(shl45_171, conv47_178) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_171, conv47_178, tmp_var);
      add48_183 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_207_inst
    process(shl54_196, conv56_203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_196, conv56_203, tmp_var);
      add57_208 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_308_inst
    process(shl96_297, conv98_304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_297, conv98_304, tmp_var);
      add99_309 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_333_inst
    process(shl105_322, conv107_329) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_322, conv107_329, tmp_var);
      add108_334 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_358_inst
    process(shl114_347, conv116_354) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_347, conv116_354, tmp_var);
      add117_359 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_383_inst
    process(shl123_372, conv125_379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_372, conv125_379, tmp_var);
      add126_384 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_408_inst
    process(shl132_397, conv134_404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_397, conv134_404, tmp_var);
      add135_409 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_57_inst
    process(shl_46, conv3_53) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_46, conv3_53, tmp_var);
      add_58 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_82_inst
    process(shl9_71, conv11_78) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_71, conv11_78, tmp_var);
      add12_83 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_508_inst
    process(shl146_497, conv149_504) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_497, conv149_504, tmp_var);
      add150_509 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_526_inst
    process(shl152_515, conv155_522) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_515, conv155_522, tmp_var);
      add156_527 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_544_inst
    process(shl158_533, conv161_540) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_533, conv161_540, tmp_var);
      add162_545 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_562_inst
    process(shl164_551, conv167_558) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_551, conv167_558, tmp_var);
      add168_563 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_580_inst
    process(shl170_569, conv173_576) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_569, conv173_576, tmp_var);
      add174_581 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_598_inst
    process(shl176_587, conv179_594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_587, conv179_594, tmp_var);
      add180_599 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_616_inst
    process(shl182_605, conv185_612) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_605, conv185_612, tmp_var);
      add186_617 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_715_inst
    process(shl202_704, conv205_711) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_704, conv205_711, tmp_var);
      add206_716 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_733_inst
    process(shl208_722, conv211_729) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_722, conv211_729, tmp_var);
      add212_734 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_751_inst
    process(shl214_740, conv217_747) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_740, conv217_747, tmp_var);
      add218_752 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_769_inst
    process(shl220_758, conv223_765) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_758, conv223_765, tmp_var);
      add224_770 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_787_inst
    process(shl226_776, conv229_783) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_776, conv229_783, tmp_var);
      add230_788 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_805_inst
    process(shl232_794, conv235_801) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_794, conv235_801, tmp_var);
      add236_806 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_823_inst
    process(shl238_812, conv241_819) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_812, conv241_819, tmp_var);
      add242_824 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_120_inst
    process(conv26_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_115, type_cast_119_wire_constant, tmp_var);
      shl27_121 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_145_inst
    process(conv35_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_140, type_cast_144_wire_constant, tmp_var);
      shl36_146 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_170_inst
    process(conv44_165) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_165, type_cast_169_wire_constant, tmp_var);
      shl45_171 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_195_inst
    process(conv53_190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_190, type_cast_194_wire_constant, tmp_var);
      shl54_196 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_296_inst
    process(conv95_291) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_291, type_cast_295_wire_constant, tmp_var);
      shl96_297 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_321_inst
    process(conv104_316) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_316, type_cast_320_wire_constant, tmp_var);
      shl105_322 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_346_inst
    process(conv113_341) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_341, type_cast_345_wire_constant, tmp_var);
      shl114_347 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_371_inst
    process(conv122_366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_366, type_cast_370_wire_constant, tmp_var);
      shl123_372 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_396_inst
    process(conv131_391) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_391, type_cast_395_wire_constant, tmp_var);
      shl132_397 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_45_inst
    process(conv1_40) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_40, type_cast_44_wire_constant, tmp_var);
      shl_46 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_70_inst
    process(conv8_65) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_65, type_cast_69_wire_constant, tmp_var);
      shl9_71 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_95_inst
    process(conv17_90) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_90, type_cast_94_wire_constant, tmp_var);
      shl18_96 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_496_inst
    process(conv144_491) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_491, type_cast_495_wire_constant, tmp_var);
      shl146_497 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_514_inst
    process(add150_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_509, type_cast_513_wire_constant, tmp_var);
      shl152_515 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_532_inst
    process(add156_527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_527, type_cast_531_wire_constant, tmp_var);
      shl158_533 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_550_inst
    process(add162_545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_545, type_cast_549_wire_constant, tmp_var);
      shl164_551 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_568_inst
    process(add168_563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_563, type_cast_567_wire_constant, tmp_var);
      shl170_569 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_586_inst
    process(add174_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_581, type_cast_585_wire_constant, tmp_var);
      shl176_587 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_604_inst
    process(add180_599) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_599, type_cast_603_wire_constant, tmp_var);
      shl182_605 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_703_inst
    process(conv200_698) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_698, type_cast_702_wire_constant, tmp_var);
      shl202_704 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_721_inst
    process(add206_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_716, type_cast_720_wire_constant, tmp_var);
      shl208_722 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_739_inst
    process(add212_734) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_734, type_cast_738_wire_constant, tmp_var);
      shl214_740 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_757_inst
    process(add218_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_752, type_cast_756_wire_constant, tmp_var);
      shl220_758 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_775_inst
    process(add224_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_770, type_cast_774_wire_constant, tmp_var);
      shl226_776 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_793_inst
    process(add230_788) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_788, type_cast_792_wire_constant, tmp_var);
      shl232_794 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_811_inst
    process(add236_806) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_806, type_cast_810_wire_constant, tmp_var);
      shl238_812 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1205_inst
    process(conv355_1201, conv276_969) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1201, conv276_969, tmp_var);
      sub_1206 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1228_inst
    process(tmp458_1223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp458_1223, type_cast_1227_wire_constant, tmp_var);
      tmp459_1229 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_414_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_230, type_cast_413_wire_constant, tmp_var);
      cmp451_416 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_430_inst
    process(mul91_284) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_284, type_cast_429_wire_constant, tmp_var);
      cmp194447_431 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_443_inst
    process(shr_236) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_236, type_cast_442_wire_constant, tmp_var);
      tmp501_444 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_650_inst
    process(tmp486_645) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp486_645, type_cast_649_wire_constant, tmp_var);
      tmp487_651 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_875_inst
    process(mul259_870) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_870, type_cast_874_wire_constant, tmp_var);
      cmp264443_876 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_894_inst
    process(tmp470_889) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp470_889, type_cast_893_wire_constant, tmp_var);
      tmp471_895 <= tmp_var; --
    end process;
    -- shared split operator group (100) : array_obj_ref_1267_index_offset 
    ApIntAdd_group_100: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1266_scaled;
      array_obj_ref_1267_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1267_index_offset_req_0;
      array_obj_ref_1267_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1267_index_offset_req_1;
      array_obj_ref_1267_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_100_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_100_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_100",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 100
    -- shared split operator group (101) : array_obj_ref_482_index_offset 
    ApIntAdd_group_101: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar493_481_scaled;
      array_obj_ref_482_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_482_index_offset_req_0;
      array_obj_ref_482_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_482_index_offset_req_1;
      array_obj_ref_482_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_101_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_101_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_101",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 101
    -- shared split operator group (102) : array_obj_ref_689_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar477_688_scaled;
      array_obj_ref_689_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_689_index_offset_req_0;
      array_obj_ref_689_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_689_index_offset_req_1;
      array_obj_ref_689_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : array_obj_ref_933_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar463_932_scaled;
      array_obj_ref_933_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_933_index_offset_req_0;
      array_obj_ref_933_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_933_index_offset_req_1;
      array_obj_ref_933_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- unary operator type_cast_1199_inst
    process(call354_1196) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1196, tmp_var);
      type_cast_1199_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_967_inst
    process(call275_963) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_963, tmp_var);
      type_cast_967_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1272_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1272_load_0_req_0;
      ptr_deref_1272_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1272_load_0_req_1;
      ptr_deref_1272_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1272_word_address_0;
      ptr_deref_1272_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_619_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_619_store_0_req_0;
      ptr_deref_619_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_619_store_0_req_1;
      ptr_deref_619_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_619_word_address_0;
      data_in <= ptr_deref_619_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_826_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_826_store_0_req_0;
      ptr_deref_826_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_826_store_0_req_1;
      ptr_deref_826_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_826_word_address_0;
      data_in <= ptr_deref_826_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_937_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_937_store_0_req_0;
      ptr_deref_937_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_937_store_0_req_1;
      ptr_deref_937_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_937_word_address_0;
      data_in <= ptr_deref_937_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1183_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1183_inst_req_0;
      RPIPE_Block0_done_1183_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1183_inst_req_1;
      RPIPE_Block0_done_1183_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1184 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1186_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1186_inst_req_0;
      RPIPE_Block1_done_1186_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1186_inst_req_1;
      RPIPE_Block1_done_1186_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1187 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1189_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1189_inst_req_0;
      RPIPE_Block2_done_1189_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1189_inst_req_1;
      RPIPE_Block2_done_1189_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1190 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1192_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1192_inst_req_0;
      RPIPE_Block3_done_1192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1192_inst_req_1;
      RPIPE_Block3_done_1192_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1193 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_98_inst RPIPE_ConvTranspose_input_pipe_48_inst RPIPE_ConvTranspose_input_pipe_85_inst RPIPE_ConvTranspose_input_pipe_185_inst RPIPE_ConvTranspose_input_pipe_173_inst RPIPE_ConvTranspose_input_pipe_160_inst RPIPE_ConvTranspose_input_pipe_73_inst RPIPE_ConvTranspose_input_pipe_60_inst RPIPE_ConvTranspose_input_pipe_135_inst RPIPE_ConvTranspose_input_pipe_110_inst RPIPE_ConvTranspose_input_pipe_148_inst RPIPE_ConvTranspose_input_pipe_123_inst RPIPE_ConvTranspose_input_pipe_198_inst RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_386_inst RPIPE_ConvTranspose_input_pipe_361_inst RPIPE_ConvTranspose_input_pipe_486_inst RPIPE_ConvTranspose_input_pipe_349_inst RPIPE_ConvTranspose_input_pipe_374_inst RPIPE_ConvTranspose_input_pipe_311_inst RPIPE_ConvTranspose_input_pipe_299_inst RPIPE_ConvTranspose_input_pipe_399_inst RPIPE_ConvTranspose_input_pipe_336_inst RPIPE_ConvTranspose_input_pipe_324_inst RPIPE_ConvTranspose_input_pipe_286_inst RPIPE_ConvTranspose_input_pipe_499_inst RPIPE_ConvTranspose_input_pipe_517_inst RPIPE_ConvTranspose_input_pipe_535_inst RPIPE_ConvTranspose_input_pipe_553_inst RPIPE_ConvTranspose_input_pipe_571_inst RPIPE_ConvTranspose_input_pipe_589_inst RPIPE_ConvTranspose_input_pipe_607_inst RPIPE_ConvTranspose_input_pipe_693_inst RPIPE_ConvTranspose_input_pipe_706_inst RPIPE_ConvTranspose_input_pipe_724_inst RPIPE_ConvTranspose_input_pipe_742_inst RPIPE_ConvTranspose_input_pipe_760_inst RPIPE_ConvTranspose_input_pipe_778_inst RPIPE_ConvTranspose_input_pipe_796_inst RPIPE_ConvTranspose_input_pipe_814_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_386_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_361_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_486_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_349_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_374_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_311_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_299_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_399_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_324_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_286_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_517_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_535_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_553_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_571_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_589_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_607_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_693_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_706_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_724_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_742_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_814_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_386_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_361_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_486_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_349_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_374_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_311_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_299_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_399_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_324_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_286_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_517_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_535_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_553_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_571_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_589_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_607_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_693_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_706_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_724_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_742_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_814_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_386_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_361_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_486_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_349_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_374_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_311_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_299_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_399_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_336_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_324_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_286_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_517_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_535_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_553_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_571_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_589_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_607_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_693_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_706_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_724_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_742_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_814_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_386_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_361_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_486_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_349_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_374_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_311_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_299_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_399_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_336_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_324_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_286_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_517_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_535_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_553_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_571_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_589_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_607_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_693_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_706_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_724_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_742_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_814_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call19_99 <= data_out(319 downto 312);
      call2_49 <= data_out(311 downto 304);
      call14_86 <= data_out(303 downto 296);
      call50_186 <= data_out(295 downto 288);
      call46_174 <= data_out(287 downto 280);
      call41_161 <= data_out(279 downto 272);
      call10_74 <= data_out(271 downto 264);
      call5_61 <= data_out(263 downto 256);
      call32_136 <= data_out(255 downto 248);
      call23_111 <= data_out(247 downto 240);
      call37_149 <= data_out(239 downto 232);
      call28_124 <= data_out(231 downto 224);
      call55_199 <= data_out(223 downto 216);
      call_36 <= data_out(215 downto 208);
      call128_387 <= data_out(207 downto 200);
      call119_362 <= data_out(199 downto 192);
      call143_487 <= data_out(191 downto 184);
      call115_350 <= data_out(183 downto 176);
      call124_375 <= data_out(175 downto 168);
      call101_312 <= data_out(167 downto 160);
      call97_300 <= data_out(159 downto 152);
      call133_400 <= data_out(151 downto 144);
      call110_337 <= data_out(143 downto 136);
      call106_325 <= data_out(135 downto 128);
      call92_287 <= data_out(127 downto 120);
      call147_500 <= data_out(119 downto 112);
      call153_518 <= data_out(111 downto 104);
      call159_536 <= data_out(103 downto 96);
      call165_554 <= data_out(95 downto 88);
      call171_572 <= data_out(87 downto 80);
      call177_590 <= data_out(79 downto 72);
      call183_608 <= data_out(71 downto 64);
      call199_694 <= data_out(63 downto 56);
      call203_707 <= data_out(55 downto 48);
      call209_725 <= data_out(47 downto 40);
      call215_743 <= data_out(39 downto 32);
      call221_761 <= data_out(31 downto 24);
      call227_779 <= data_out(23 downto 16);
      call233_797 <= data_out(15 downto 8);
      call239_815 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_970_inst WPIPE_Block0_start_973_inst WPIPE_Block0_start_976_inst WPIPE_Block0_start_979_inst WPIPE_Block0_start_982_inst WPIPE_Block0_start_985_inst WPIPE_Block0_start_988_inst WPIPE_Block0_start_991_inst WPIPE_Block0_start_994_inst WPIPE_Block0_start_997_inst WPIPE_Block0_start_1001_inst WPIPE_Block0_start_1005_inst WPIPE_Block0_start_1008_inst WPIPE_Block0_start_1011_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_970_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_973_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_976_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_979_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_982_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_985_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_988_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_991_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_994_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_997_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_1001_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_1005_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_1008_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1011_inst_req_0;
      WPIPE_Block0_start_970_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_973_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_976_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_979_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_982_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_985_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_988_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_991_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_994_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_997_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_1001_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_1005_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_1008_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1011_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_970_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_973_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_976_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_979_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_982_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_985_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_988_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_991_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_994_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_997_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_1001_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_1005_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_1008_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1011_inst_req_1;
      WPIPE_Block0_start_970_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_973_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_976_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_979_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_982_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_985_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_988_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_991_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_994_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_997_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_1001_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_1005_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_1008_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1011_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add99_309 & add108_334 & type_cast_999_wire_constant & type_cast_1003_wire_constant & add117_359 & add126_384 & add135_409;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1014_inst WPIPE_Block1_start_1017_inst WPIPE_Block1_start_1020_inst WPIPE_Block1_start_1023_inst WPIPE_Block1_start_1026_inst WPIPE_Block1_start_1029_inst WPIPE_Block1_start_1032_inst WPIPE_Block1_start_1035_inst WPIPE_Block1_start_1038_inst WPIPE_Block1_start_1045_inst WPIPE_Block1_start_1058_inst WPIPE_Block1_start_1061_inst WPIPE_Block1_start_1064_inst WPIPE_Block1_start_1067_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1014_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1017_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1020_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1023_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1026_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1029_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1032_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1035_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1038_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1045_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1058_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1061_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1064_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1067_inst_req_0;
      WPIPE_Block1_start_1014_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1017_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1020_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1023_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1026_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1029_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1032_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1035_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1038_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1045_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1058_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1061_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1064_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1067_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1014_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1017_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1020_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1023_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1026_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1029_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1032_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1035_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1038_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1045_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1058_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1061_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1064_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1067_inst_req_1;
      WPIPE_Block1_start_1014_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1017_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1020_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1023_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1026_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1029_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1032_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1035_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1038_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1045_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1058_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1061_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1064_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1067_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add99_309 & add108_334 & conv304_1044 & conv307_1057 & add117_359 & add126_384 & add135_409;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1091_inst WPIPE_Block2_start_1117_inst WPIPE_Block2_start_1114_inst WPIPE_Block2_start_1123_inst WPIPE_Block2_start_1094_inst WPIPE_Block2_start_1101_inst WPIPE_Block2_start_1120_inst WPIPE_Block2_start_1088_inst WPIPE_Block2_start_1070_inst WPIPE_Block2_start_1073_inst WPIPE_Block2_start_1076_inst WPIPE_Block2_start_1079_inst WPIPE_Block2_start_1082_inst WPIPE_Block2_start_1085_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1091_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1117_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1114_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1123_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1094_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1101_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1120_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1088_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1070_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1073_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1076_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1079_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1082_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1085_inst_req_0;
      WPIPE_Block2_start_1091_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1117_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1114_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1123_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1094_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1101_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1120_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1088_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1070_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1073_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1076_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1079_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1082_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1085_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1091_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1117_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1114_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1123_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1094_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1101_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1120_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1088_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1070_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1073_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1076_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1079_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1082_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1085_inst_req_1;
      WPIPE_Block2_start_1091_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1117_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1114_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1123_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1094_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1101_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1120_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1088_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1070_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1073_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1076_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1079_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1082_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1085_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add99_309 & add117_359 & conv324_1113 & add135_409 & add108_334 & conv321_1100 & add126_384 & add57_208 & add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1150_inst WPIPE_Block3_start_1147_inst WPIPE_Block3_start_1129_inst WPIPE_Block3_start_1126_inst WPIPE_Block3_start_1132_inst WPIPE_Block3_start_1135_inst WPIPE_Block3_start_1157_inst WPIPE_Block3_start_1138_inst WPIPE_Block3_start_1141_inst WPIPE_Block3_start_1144_inst WPIPE_Block3_start_1170_inst WPIPE_Block3_start_1179_inst WPIPE_Block3_start_1176_inst WPIPE_Block3_start_1173_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1150_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1147_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1129_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1126_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1132_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1135_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1157_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1138_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1141_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1144_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1170_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1179_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1176_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1173_inst_req_0;
      WPIPE_Block3_start_1150_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1147_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1129_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1126_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1132_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1135_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1157_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1138_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1141_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1144_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1170_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1179_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1176_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1173_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1150_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1147_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1129_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1126_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1132_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1135_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1157_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1138_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1141_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1144_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1170_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1179_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1176_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1173_inst_req_1;
      WPIPE_Block3_start_1150_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1147_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1129_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1126_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1132_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1135_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1157_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1138_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1141_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1144_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1170_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1179_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1176_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1173_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add108_334 & add99_309 & add12_83 & add_58 & add21_108 & add30_133 & conv338_1156 & add39_158 & add48_183 & add57_208 & conv341_1169 & add135_409 & add126_384 & add117_359;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1351_inst WPIPE_ConvTranspose_output_pipe_1348_inst WPIPE_ConvTranspose_output_pipe_1354_inst WPIPE_ConvTranspose_output_pipe_1357_inst WPIPE_ConvTranspose_output_pipe_1360_inst WPIPE_ConvTranspose_output_pipe_1363_inst WPIPE_ConvTranspose_output_pipe_1366_inst WPIPE_ConvTranspose_output_pipe_1369_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1351_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1348_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1354_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1357_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1360_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1363_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1366_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1369_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1351_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1348_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1354_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1357_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1360_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1363_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1366_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1369_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1351_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1348_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1354_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1357_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1360_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1363_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1366_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1369_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1351_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1348_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1354_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1357_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1360_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1363_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1366_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1369_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv411_1337 & conv417_1347 & conv405_1327 & conv399_1317 & conv393_1307 & conv387_1297 & conv381_1287 & conv375_1277;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1207_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1207_inst_req_0;
      WPIPE_elapsed_time_pipe_1207_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1207_inst_req_1;
      WPIPE_elapsed_time_pipe_1207_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1206;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_1196_call call_stmt_963_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1196_call_req_0;
      reqL_unguarded(0) <= call_stmt_963_call_req_0;
      call_stmt_1196_call_ack_0 <= ackL_unguarded(1);
      call_stmt_963_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1196_call_req_1;
      reqR_unguarded(0) <= call_stmt_963_call_req_1;
      call_stmt_1196_call_ack_1 <= ackR_unguarded(1);
      call_stmt_963_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call354_1196 <= data_out(127 downto 64);
      call275_963 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3548_start: Boolean;
  signal convTransposeA_CP_3548_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1576_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1457_inst_req_1 : boolean;
  signal type_cast_1496_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1439_inst_ack_0 : boolean;
  signal type_cast_1443_inst_req_0 : boolean;
  signal ptr_deref_1617_load_0_ack_0 : boolean;
  signal type_cast_1484_inst_req_0 : boolean;
  signal type_cast_1492_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1457_inst_ack_1 : boolean;
  signal type_cast_1576_inst_req_0 : boolean;
  signal array_obj_ref_1612_index_offset_req_1 : boolean;
  signal array_obj_ref_1635_index_offset_ack_0 : boolean;
  signal type_cast_1606_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1454_inst_req_1 : boolean;
  signal type_cast_1443_inst_ack_0 : boolean;
  signal type_cast_1496_inst_req_1 : boolean;
  signal type_cast_1492_inst_ack_1 : boolean;
  signal ptr_deref_1617_load_0_req_0 : boolean;
  signal RPIPE_Block0_start_1457_inst_req_0 : boolean;
  signal array_obj_ref_1612_index_offset_ack_1 : boolean;
  signal RPIPE_Block0_start_1454_inst_ack_1 : boolean;
  signal type_cast_1488_inst_req_0 : boolean;
  signal type_cast_1572_inst_ack_0 : boolean;
  signal type_cast_1576_inst_req_1 : boolean;
  signal type_cast_1568_inst_ack_1 : boolean;
  signal type_cast_1488_inst_ack_1 : boolean;
  signal addr_of_1636_final_reg_ack_1 : boolean;
  signal type_cast_1568_inst_req_1 : boolean;
  signal array_obj_ref_1635_index_offset_req_1 : boolean;
  signal type_cast_1492_inst_ack_0 : boolean;
  signal type_cast_1484_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1439_inst_req_0 : boolean;
  signal type_cast_1572_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1439_inst_req_1 : boolean;
  signal addr_of_1636_final_reg_ack_0 : boolean;
  signal array_obj_ref_1635_index_offset_ack_1 : boolean;
  signal type_cast_1484_inst_req_1 : boolean;
  signal type_cast_1572_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1454_inst_ack_0 : boolean;
  signal type_cast_1576_inst_ack_1 : boolean;
  signal type_cast_1606_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1454_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1451_inst_req_1 : boolean;
  signal addr_of_1636_final_reg_req_0 : boolean;
  signal type_cast_1568_inst_req_0 : boolean;
  signal array_obj_ref_1635_index_offset_req_0 : boolean;
  signal addr_of_1613_final_reg_req_0 : boolean;
  signal type_cast_1488_inst_req_1 : boolean;
  signal type_cast_1568_inst_ack_0 : boolean;
  signal type_cast_1606_inst_req_1 : boolean;
  signal type_cast_1430_inst_req_1 : boolean;
  signal addr_of_1636_final_reg_req_1 : boolean;
  signal addr_of_1613_final_reg_req_1 : boolean;
  signal array_obj_ref_1612_index_offset_req_0 : boolean;
  signal type_cast_1492_inst_req_0 : boolean;
  signal type_cast_1430_inst_ack_1 : boolean;
  signal array_obj_ref_1612_index_offset_ack_0 : boolean;
  signal type_cast_1606_inst_ack_1 : boolean;
  signal type_cast_1443_inst_req_1 : boolean;
  signal type_cast_1572_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1457_inst_ack_0 : boolean;
  signal type_cast_1496_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1439_inst_ack_1 : boolean;
  signal type_cast_1496_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1451_inst_ack_1 : boolean;
  signal type_cast_1443_inst_ack_1 : boolean;
  signal addr_of_1613_final_reg_ack_1 : boolean;
  signal RPIPE_Block0_start_1451_inst_ack_0 : boolean;
  signal ptr_deref_1617_load_0_ack_1 : boolean;
  signal type_cast_1488_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1451_inst_req_0 : boolean;
  signal addr_of_1613_final_reg_ack_0 : boolean;
  signal type_cast_1484_inst_ack_0 : boolean;
  signal ptr_deref_1617_load_0_req_1 : boolean;
  signal RPIPE_Block0_start_1399_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1399_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1399_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1399_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1402_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1402_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1402_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1402_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1405_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1405_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1405_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1405_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1408_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1408_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1408_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1408_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1411_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1411_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1411_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1411_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1414_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1414_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1414_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1414_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1417_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1417_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1417_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1417_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1420_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1420_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1420_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1420_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1423_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1423_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1423_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1423_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1426_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1426_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1426_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1426_inst_ack_1 : boolean;
  signal type_cast_1430_inst_req_0 : boolean;
  signal type_cast_1430_inst_ack_0 : boolean;
  signal ptr_deref_1639_store_0_req_0 : boolean;
  signal ptr_deref_1639_store_0_ack_0 : boolean;
  signal ptr_deref_1639_store_0_req_1 : boolean;
  signal ptr_deref_1639_store_0_ack_1 : boolean;
  signal type_cast_1644_inst_req_0 : boolean;
  signal type_cast_1644_inst_ack_0 : boolean;
  signal type_cast_1644_inst_req_1 : boolean;
  signal type_cast_1644_inst_ack_1 : boolean;
  signal if_stmt_1657_branch_req_0 : boolean;
  signal if_stmt_1657_branch_ack_1 : boolean;
  signal if_stmt_1657_branch_ack_0 : boolean;
  signal type_cast_1685_inst_req_0 : boolean;
  signal type_cast_1685_inst_ack_0 : boolean;
  signal type_cast_1685_inst_req_1 : boolean;
  signal type_cast_1685_inst_ack_1 : boolean;
  signal type_cast_1701_inst_req_0 : boolean;
  signal type_cast_1701_inst_ack_0 : boolean;
  signal type_cast_1701_inst_req_1 : boolean;
  signal type_cast_1701_inst_ack_1 : boolean;
  signal if_stmt_1708_branch_req_0 : boolean;
  signal if_stmt_1708_branch_ack_1 : boolean;
  signal if_stmt_1708_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1744_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1744_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1744_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1744_inst_ack_1 : boolean;
  signal phi_stmt_1506_req_0 : boolean;
  signal phi_stmt_1513_req_0 : boolean;
  signal phi_stmt_1520_req_0 : boolean;
  signal phi_stmt_1527_req_0 : boolean;
  signal type_cast_1512_inst_req_0 : boolean;
  signal type_cast_1512_inst_ack_0 : boolean;
  signal type_cast_1512_inst_req_1 : boolean;
  signal type_cast_1512_inst_ack_1 : boolean;
  signal phi_stmt_1506_req_1 : boolean;
  signal type_cast_1519_inst_req_0 : boolean;
  signal type_cast_1519_inst_ack_0 : boolean;
  signal type_cast_1519_inst_req_1 : boolean;
  signal type_cast_1519_inst_ack_1 : boolean;
  signal phi_stmt_1513_req_1 : boolean;
  signal type_cast_1526_inst_req_0 : boolean;
  signal type_cast_1526_inst_ack_0 : boolean;
  signal type_cast_1526_inst_req_1 : boolean;
  signal type_cast_1526_inst_ack_1 : boolean;
  signal phi_stmt_1520_req_1 : boolean;
  signal type_cast_1533_inst_req_0 : boolean;
  signal type_cast_1533_inst_ack_0 : boolean;
  signal type_cast_1533_inst_req_1 : boolean;
  signal type_cast_1533_inst_ack_1 : boolean;
  signal phi_stmt_1527_req_1 : boolean;
  signal phi_stmt_1506_ack_0 : boolean;
  signal phi_stmt_1513_ack_0 : boolean;
  signal phi_stmt_1520_ack_0 : boolean;
  signal phi_stmt_1527_ack_0 : boolean;
  signal phi_stmt_1715_req_1 : boolean;
  signal type_cast_1725_inst_req_0 : boolean;
  signal type_cast_1725_inst_ack_0 : boolean;
  signal type_cast_1725_inst_req_1 : boolean;
  signal type_cast_1725_inst_ack_1 : boolean;
  signal phi_stmt_1722_req_0 : boolean;
  signal type_cast_1733_inst_req_0 : boolean;
  signal type_cast_1733_inst_ack_0 : boolean;
  signal type_cast_1733_inst_req_1 : boolean;
  signal type_cast_1733_inst_ack_1 : boolean;
  signal phi_stmt_1728_req_1 : boolean;
  signal type_cast_1718_inst_req_0 : boolean;
  signal type_cast_1718_inst_ack_0 : boolean;
  signal type_cast_1718_inst_req_1 : boolean;
  signal type_cast_1718_inst_ack_1 : boolean;
  signal phi_stmt_1715_req_0 : boolean;
  signal type_cast_1727_inst_req_0 : boolean;
  signal type_cast_1727_inst_ack_0 : boolean;
  signal type_cast_1727_inst_req_1 : boolean;
  signal type_cast_1727_inst_ack_1 : boolean;
  signal phi_stmt_1722_req_1 : boolean;
  signal type_cast_1731_inst_req_0 : boolean;
  signal type_cast_1731_inst_ack_0 : boolean;
  signal type_cast_1731_inst_req_1 : boolean;
  signal type_cast_1731_inst_ack_1 : boolean;
  signal phi_stmt_1728_req_0 : boolean;
  signal phi_stmt_1715_ack_0 : boolean;
  signal phi_stmt_1722_ack_0 : boolean;
  signal phi_stmt_1728_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3548_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3548_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3548_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3548_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3548: Block -- control-path 
    signal convTransposeA_CP_3548_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3548_elements(0) <= convTransposeA_CP_3548_start;
    convTransposeA_CP_3548_symbol <= convTransposeA_CP_3548_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1397/$entry
      -- CP-element group 0: 	 branch_block_stmt_1397/branch_block_stmt_1397__entry__
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458__entry__
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/$entry
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_update_start_
      -- 
    cr_3741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(0), ack => type_cast_1430_inst_req_1); -- 
    cr_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(0), ack => type_cast_1443_inst_req_1); -- 
    rr_3596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(0), ack => RPIPE_Block0_start_1399_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1397/merge_stmt_1714__exit__
      -- CP-element group 1: 	 branch_block_stmt_1397/assign_stmt_1740__entry__
      -- CP-element group 1: 	 branch_block_stmt_1397/assign_stmt_1740__exit__
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1397/assign_stmt_1740/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/assign_stmt_1740/$exit
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Update/cr
      -- 
    rr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1512_inst_req_0); -- 
    cr_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1512_inst_req_1); -- 
    rr_4305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1519_inst_req_0); -- 
    cr_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1519_inst_req_1); -- 
    rr_4328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1526_inst_req_0); -- 
    cr_4333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1526_inst_req_1); -- 
    rr_4351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1533_inst_req_0); -- 
    cr_4356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(1), ack => type_cast_1533_inst_req_1); -- 
    convTransposeA_CP_3548_elements(1) <= convTransposeA_CP_3548_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Update/cr
      -- 
    ra_3597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1399_inst_ack_0, ack => convTransposeA_CP_3548_elements(2)); -- 
    cr_3601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(2), ack => RPIPE_Block0_start_1399_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1399_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Sample/rr
      -- 
    ca_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1399_inst_ack_1, ack => convTransposeA_CP_3548_elements(3)); -- 
    rr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(3), ack => RPIPE_Block0_start_1402_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Update/cr
      -- 
    ra_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1402_inst_ack_0, ack => convTransposeA_CP_3548_elements(4)); -- 
    cr_3615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(4), ack => RPIPE_Block0_start_1402_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1402_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Sample/rr
      -- 
    ca_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1402_inst_ack_1, ack => convTransposeA_CP_3548_elements(5)); -- 
    rr_3624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(5), ack => RPIPE_Block0_start_1405_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Update/cr
      -- 
    ra_3625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1405_inst_ack_0, ack => convTransposeA_CP_3548_elements(6)); -- 
    cr_3629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(6), ack => RPIPE_Block0_start_1405_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1405_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Sample/rr
      -- 
    ca_3630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1405_inst_ack_1, ack => convTransposeA_CP_3548_elements(7)); -- 
    rr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(7), ack => RPIPE_Block0_start_1408_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Update/cr
      -- 
    ra_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1408_inst_ack_0, ack => convTransposeA_CP_3548_elements(8)); -- 
    cr_3643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(8), ack => RPIPE_Block0_start_1408_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1408_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Sample/rr
      -- 
    ca_3644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1408_inst_ack_1, ack => convTransposeA_CP_3548_elements(9)); -- 
    rr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(9), ack => RPIPE_Block0_start_1411_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Update/cr
      -- 
    ra_3653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1411_inst_ack_0, ack => convTransposeA_CP_3548_elements(10)); -- 
    cr_3657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(10), ack => RPIPE_Block0_start_1411_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1411_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Sample/rr
      -- 
    ca_3658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1411_inst_ack_1, ack => convTransposeA_CP_3548_elements(11)); -- 
    rr_3666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(11), ack => RPIPE_Block0_start_1414_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Update/cr
      -- 
    ra_3667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1414_inst_ack_0, ack => convTransposeA_CP_3548_elements(12)); -- 
    cr_3671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(12), ack => RPIPE_Block0_start_1414_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1414_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Sample/rr
      -- 
    ca_3672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1414_inst_ack_1, ack => convTransposeA_CP_3548_elements(13)); -- 
    rr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(13), ack => RPIPE_Block0_start_1417_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Update/cr
      -- 
    ra_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1417_inst_ack_0, ack => convTransposeA_CP_3548_elements(14)); -- 
    cr_3685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(14), ack => RPIPE_Block0_start_1417_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1417_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Sample/rr
      -- 
    ca_3686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1417_inst_ack_1, ack => convTransposeA_CP_3548_elements(15)); -- 
    rr_3694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(15), ack => RPIPE_Block0_start_1420_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Update/cr
      -- 
    ra_3695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1420_inst_ack_0, ack => convTransposeA_CP_3548_elements(16)); -- 
    cr_3699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(16), ack => RPIPE_Block0_start_1420_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1420_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Sample/rr
      -- 
    ca_3700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1420_inst_ack_1, ack => convTransposeA_CP_3548_elements(17)); -- 
    rr_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(17), ack => RPIPE_Block0_start_1423_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Update/cr
      -- 
    ra_3709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1423_inst_ack_0, ack => convTransposeA_CP_3548_elements(18)); -- 
    cr_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(18), ack => RPIPE_Block0_start_1423_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1423_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Sample/rr
      -- 
    ca_3714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1423_inst_ack_1, ack => convTransposeA_CP_3548_elements(19)); -- 
    rr_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(19), ack => RPIPE_Block0_start_1426_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Update/cr
      -- 
    ra_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1426_inst_ack_0, ack => convTransposeA_CP_3548_elements(20)); -- 
    cr_3727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(20), ack => RPIPE_Block0_start_1426_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1426_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Sample/rr
      -- 
    ca_3728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1426_inst_ack_1, ack => convTransposeA_CP_3548_elements(21)); -- 
    rr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(21), ack => type_cast_1430_inst_req_0); -- 
    rr_3750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(21), ack => RPIPE_Block0_start_1439_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Sample/ra
      -- 
    ra_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_0, ack => convTransposeA_CP_3548_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1430_update_completed_
      -- 
    ca_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_1, ack => convTransposeA_CP_3548_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_update_start_
      -- 
    ra_3751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1439_inst_ack_0, ack => convTransposeA_CP_3548_elements(24)); -- 
    cr_3755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(24), ack => RPIPE_Block0_start_1439_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1439_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Sample/rr
      -- 
    ca_3756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1439_inst_ack_1, ack => convTransposeA_CP_3548_elements(25)); -- 
    rr_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(25), ack => type_cast_1443_inst_req_0); -- 
    rr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(25), ack => RPIPE_Block0_start_1451_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_sample_completed_
      -- 
    ra_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1443_inst_ack_0, ack => convTransposeA_CP_3548_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/type_cast_1443_Update/ca
      -- 
    ca_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1443_inst_ack_1, ack => convTransposeA_CP_3548_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Sample/ra
      -- 
    ra_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1451_inst_ack_0, ack => convTransposeA_CP_3548_elements(28)); -- 
    cr_3783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(28), ack => RPIPE_Block0_start_1451_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1451_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Sample/$entry
      -- 
    ca_3784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1451_inst_ack_1, ack => convTransposeA_CP_3548_elements(29)); -- 
    rr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(29), ack => RPIPE_Block0_start_1454_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Sample/$exit
      -- 
    ra_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1454_inst_ack_0, ack => convTransposeA_CP_3548_elements(30)); -- 
    cr_3797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(30), ack => RPIPE_Block0_start_1454_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1454_update_completed_
      -- 
    ca_3798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1454_inst_ack_1, ack => convTransposeA_CP_3548_elements(31)); -- 
    rr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(31), ack => RPIPE_Block0_start_1457_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Sample/ra
      -- 
    ra_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1457_inst_ack_0, ack => convTransposeA_CP_3548_elements(32)); -- 
    cr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(32), ack => RPIPE_Block0_start_1457_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/RPIPE_Block0_start_1457_update_completed_
      -- 
    ca_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1457_inst_ack_1, ack => convTransposeA_CP_3548_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458__exit__
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503__entry__
      -- CP-element group 34: 	 branch_block_stmt_1397/assign_stmt_1400_to_assign_stmt_1458/$exit
      -- 
    rr_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1484_inst_req_0); -- 
    cr_3856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1492_inst_req_1); -- 
    cr_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1496_inst_req_1); -- 
    rr_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1488_inst_req_0); -- 
    cr_3828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1484_inst_req_1); -- 
    cr_3842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1488_inst_req_1); -- 
    rr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1492_inst_req_0); -- 
    rr_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(34), ack => type_cast_1496_inst_req_0); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(23) & convTransposeA_CP_3548_elements(27) & convTransposeA_CP_3548_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Sample/ra
      -- 
    ra_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1484_inst_ack_0, ack => convTransposeA_CP_3548_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1484_Update/$exit
      -- 
    ca_3829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1484_inst_ack_1, ack => convTransposeA_CP_3548_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Sample/ra
      -- 
    ra_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_0, ack => convTransposeA_CP_3548_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1488_Update/$exit
      -- 
    ca_3843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_1, ack => convTransposeA_CP_3548_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Sample/$exit
      -- 
    ra_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1492_inst_ack_0, ack => convTransposeA_CP_3548_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1492_update_completed_
      -- 
    ca_3857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1492_inst_ack_1, ack => convTransposeA_CP_3548_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_sample_completed_
      -- 
    ra_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1496_inst_ack_0, ack => convTransposeA_CP_3548_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/type_cast_1496_update_completed_
      -- 
    ca_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1496_inst_ack_1, ack => convTransposeA_CP_3548_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503/$exit
      -- CP-element group 43: 	 branch_block_stmt_1397/assign_stmt_1465_to_assign_stmt_1503__exit__
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1506/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1513/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1520/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1527/$entry
      -- CP-element group 43: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(36) & convTransposeA_CP_3548_elements(38) & convTransposeA_CP_3548_elements(40) & convTransposeA_CP_3548_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Sample/ra
      -- 
    ra_3883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1568_inst_ack_0, ack => convTransposeA_CP_3548_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Update/ca
      -- 
    ca_3888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1568_inst_ack_1, ack => convTransposeA_CP_3548_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_sample_completed_
      -- 
    ra_3897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1572_inst_ack_0, ack => convTransposeA_CP_3548_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Update/ca
      -- 
    ca_3902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1572_inst_ack_1, ack => convTransposeA_CP_3548_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Sample/$exit
      -- 
    ra_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1576_inst_ack_0, ack => convTransposeA_CP_3548_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_update_completed_
      -- 
    ca_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1576_inst_ack_1, ack => convTransposeA_CP_3548_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Sample/$exit
      -- 
    ra_3925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_0, ack => convTransposeA_CP_3548_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_index_resized_1
      -- 
    ca_3930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_1, ack => convTransposeA_CP_3548_elements(51)); -- 
    req_3955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(51), ack => array_obj_ref_1612_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Sample/ack
      -- 
    ack_3956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1612_index_offset_ack_0, ack => convTransposeA_CP_3548_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_request/req
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_base_plus_offset/$entry
      -- 
    ack_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1612_index_offset_ack_1, ack => convTransposeA_CP_3548_elements(53)); -- 
    req_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(53), ack => addr_of_1613_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_request/ack
      -- 
    ack_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1613_final_reg_ack_0, ack => convTransposeA_CP_3548_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/word_access_start/word_0/rr
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_base_plus_offset/sum_rename_ack
      -- 
    ack_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1613_final_reg_ack_1, ack => convTransposeA_CP_3548_elements(55)); -- 
    rr_4009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(55), ack => ptr_deref_1617_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/word_access_start/word_0/ra
      -- CP-element group 56: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_sample_completed_
      -- 
    ra_4010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1617_load_0_ack_0, ack => convTransposeA_CP_3548_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/ptr_deref_1617_Merge/merge_ack
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/ptr_deref_1617_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/ptr_deref_1617_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/ptr_deref_1617_Merge/$entry
      -- 
    ca_4021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1617_load_0_ack_1, ack => convTransposeA_CP_3548_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_index_resized_1
      -- 
    req_4051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(58), ack => array_obj_ref_1635_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(45) & convTransposeA_CP_3548_elements(47) & convTransposeA_CP_3548_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_sample_complete
      -- 
    ack_4052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1635_index_offset_ack_0, ack => convTransposeA_CP_3548_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_request/req
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_base_plus_offset/$exit
      -- 
    ack_4057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1635_index_offset_ack_1, ack => convTransposeA_CP_3548_elements(60)); -- 
    req_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(60), ack => addr_of_1636_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_request/ack
      -- CP-element group 61: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_sample_completed_
      -- 
    ack_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1636_final_reg_ack_0, ack => convTransposeA_CP_3548_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_base_plus_offset/$exit
      -- 
    ack_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1636_final_reg_ack_1, ack => convTransposeA_CP_3548_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/ptr_deref_1639_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/ptr_deref_1639_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/ptr_deref_1639_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/ptr_deref_1639_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/word_access_start/word_0/rr
      -- 
    rr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(63), ack => ptr_deref_1639_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(57) & convTransposeA_CP_3548_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Sample/word_access_start/word_0/ra
      -- 
    ra_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1639_store_0_ack_0, ack => convTransposeA_CP_3548_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/word_access_complete/word_0/ca
      -- 
    ca_4122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1639_store_0_ack_1, ack => convTransposeA_CP_3548_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Sample/ra
      -- 
    ra_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_0, ack => convTransposeA_CP_3548_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Update/ca
      -- 
    ca_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_1, ack => convTransposeA_CP_3548_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1397/R_cmp_1658_place
      -- CP-element group 68: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/$exit
      -- CP-element group 68: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656__exit__
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657__entry__
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1397/if_stmt_1657_else_link/$entry
      -- 
    branch_req_4144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(68), ack => if_stmt_1657_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(52) & convTransposeA_CP_3548_elements(59) & convTransposeA_CP_3548_elements(65) & convTransposeA_CP_3548_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1397/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1397/merge_stmt_1663__exit__
      -- CP-element group 69: 	 branch_block_stmt_1397/assign_stmt_1669__entry__
      -- CP-element group 69: 	 branch_block_stmt_1397/assign_stmt_1669__exit__
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1397/if_stmt_1657_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1397/if_stmt_1657_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1397/assign_stmt_1669/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/assign_stmt_1669/$exit
      -- CP-element group 69: 	 branch_block_stmt_1397/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1397/merge_stmt_1663_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1397/merge_stmt_1663_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/merge_stmt_1663_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1397/merge_stmt_1663_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1657_branch_ack_1, ack => convTransposeA_CP_3548_elements(69)); -- 
    rr_4466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(69), ack => type_cast_1718_inst_req_0); -- 
    cr_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(69), ack => type_cast_1718_inst_req_1); -- 
    rr_4489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(69), ack => type_cast_1727_inst_req_0); -- 
    cr_4494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(69), ack => type_cast_1727_inst_req_1); -- 
    rr_4512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(69), ack => type_cast_1731_inst_req_0); -- 
    cr_4517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(69), ack => type_cast_1731_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1397/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1397/merge_stmt_1671__exit__
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707__entry__
      -- CP-element group 70: 	 branch_block_stmt_1397/if_stmt_1657_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1397/if_stmt_1657_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/$entry
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1397/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1397/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1397/merge_stmt_1671_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1397/merge_stmt_1671_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1397/merge_stmt_1671_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1397/merge_stmt_1671_PhiAck/dummy
      -- 
    else_choice_transition_4153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1657_branch_ack_0, ack => convTransposeA_CP_3548_elements(70)); -- 
    rr_4169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(70), ack => type_cast_1685_inst_req_0); -- 
    cr_4174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(70), ack => type_cast_1685_inst_req_1); -- 
    cr_4188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(70), ack => type_cast_1701_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Sample/ra
      -- 
    ra_4170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1685_inst_ack_0, ack => convTransposeA_CP_3548_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1685_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Sample/rr
      -- 
    ca_4175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1685_inst_ack_1, ack => convTransposeA_CP_3548_elements(72)); -- 
    rr_4183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(72), ack => type_cast_1701_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Sample/ra
      -- 
    ra_4184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_0, ack => convTransposeA_CP_3548_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1397/R_cmp112_1709_place
      -- CP-element group 74: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707__exit__
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708__entry__
      -- CP-element group 74: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/$exit
      -- CP-element group 74: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1397/assign_stmt_1677_to_assign_stmt_1707/type_cast_1701_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1397/if_stmt_1708_else_link/$entry
      -- 
    ca_4189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_1, ack => convTransposeA_CP_3548_elements(74)); -- 
    branch_req_4197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(74), ack => if_stmt_1708_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1397/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1397/merge_stmt_1742__exit__
      -- CP-element group 75: 	 branch_block_stmt_1397/assign_stmt_1747__entry__
      -- CP-element group 75: 	 branch_block_stmt_1397/if_stmt_1708_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1397/if_stmt_1708_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1397/assign_stmt_1747/$entry
      -- CP-element group 75: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1397/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1397/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1397/merge_stmt_1742_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1397/merge_stmt_1742_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1397/merge_stmt_1742_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1397/merge_stmt_1742_PhiAck/dummy
      -- 
    if_choice_transition_4202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1708_branch_ack_1, ack => convTransposeA_CP_3548_elements(75)); -- 
    req_4222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(75), ack => WPIPE_Block0_done_1744_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	108 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123
      -- CP-element group 76: 	 branch_block_stmt_1397/if_stmt_1708_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1397/if_stmt_1708_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1715/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1708_branch_ack_0, ack => convTransposeA_CP_3548_elements(76)); -- 
    rr_4417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(76), ack => type_cast_1725_inst_req_0); -- 
    cr_4422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(76), ack => type_cast_1725_inst_req_1); -- 
    rr_4440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(76), ack => type_cast_1733_inst_req_0); -- 
    cr_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(76), ack => type_cast_1733_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Update/req
      -- 
    ack_4223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1744_inst_ack_0, ack => convTransposeA_CP_3548_elements(77)); -- 
    req_4227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(77), ack => WPIPE_Block0_done_1744_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1397/$exit
      -- CP-element group 78: 	 branch_block_stmt_1397/branch_block_stmt_1397__exit__
      -- CP-element group 78: 	 branch_block_stmt_1397/assign_stmt_1747__exit__
      -- CP-element group 78: 	 branch_block_stmt_1397/return__
      -- CP-element group 78: 	 branch_block_stmt_1397/merge_stmt_1749__exit__
      -- CP-element group 78: 	 branch_block_stmt_1397/assign_stmt_1747/$exit
      -- CP-element group 78: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1397/assign_stmt_1747/WPIPE_Block0_done_1744_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1397/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1397/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1397/merge_stmt_1749_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1397/merge_stmt_1749_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1397/merge_stmt_1749_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1397/merge_stmt_1749_PhiAck/dummy
      -- 
    ack_4228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1744_inst_ack_1, ack => convTransposeA_CP_3548_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1506/$exit
      -- CP-element group 79: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1510_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_req
      -- 
    phi_stmt_1506_req_4239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1506_req_4239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(79), ack => phi_stmt_1506_req_0); -- 
    -- Element group convTransposeA_CP_3548_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3548_elements(43), ack => convTransposeA_CP_3548_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1513/$exit
      -- CP-element group 80: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1517_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_req
      -- 
    phi_stmt_1513_req_4247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1513_req_4247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(80), ack => phi_stmt_1513_req_0); -- 
    -- Element group convTransposeA_CP_3548_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3548_elements(43), ack => convTransposeA_CP_3548_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1520/$exit
      -- CP-element group 81: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1524_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_req
      -- 
    phi_stmt_1520_req_4255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1520_req_4255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(81), ack => phi_stmt_1520_req_0); -- 
    -- Element group convTransposeA_CP_3548_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3548_elements(43), ack => convTransposeA_CP_3548_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1527/$exit
      -- CP-element group 82: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1531_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_req
      -- 
    phi_stmt_1527_req_4263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1527_req_4263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(82), ack => phi_stmt_1527_req_0); -- 
    -- Element group convTransposeA_CP_3548_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3548_elements(43), ack => convTransposeA_CP_3548_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1397/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(79) & convTransposeA_CP_3548_elements(80) & convTransposeA_CP_3548_elements(81) & convTransposeA_CP_3548_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Sample/ra
      -- 
    ra_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1512_inst_ack_0, ack => convTransposeA_CP_3548_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/Update/ca
      -- 
    ca_4288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1512_inst_ack_1, ack => convTransposeA_CP_3548_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/$exit
      -- CP-element group 86: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/$exit
      -- CP-element group 86: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_sources/type_cast_1512/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1506/phi_stmt_1506_req
      -- 
    phi_stmt_1506_req_4289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1506_req_4289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(86), ack => phi_stmt_1506_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(84) & convTransposeA_CP_3548_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Sample/ra
      -- 
    ra_4306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1519_inst_ack_0, ack => convTransposeA_CP_3548_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/Update/ca
      -- 
    ca_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1519_inst_ack_1, ack => convTransposeA_CP_3548_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/$exit
      -- CP-element group 89: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/$exit
      -- CP-element group 89: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_sources/type_cast_1519/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1513/phi_stmt_1513_req
      -- 
    phi_stmt_1513_req_4312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1513_req_4312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(89), ack => phi_stmt_1513_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(87) & convTransposeA_CP_3548_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Sample/ra
      -- 
    ra_4329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_0, ack => convTransposeA_CP_3548_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/Update/ca
      -- 
    ca_4334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_1, ack => convTransposeA_CP_3548_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/$exit
      -- CP-element group 92: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/$exit
      -- CP-element group 92: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1526/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1520/phi_stmt_1520_req
      -- 
    phi_stmt_1520_req_4335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1520_req_4335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(92), ack => phi_stmt_1520_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(90) & convTransposeA_CP_3548_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Sample/ra
      -- 
    ra_4352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1533_inst_ack_0, ack => convTransposeA_CP_3548_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/Update/ca
      -- 
    ca_4357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1533_inst_ack_1, ack => convTransposeA_CP_3548_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/$exit
      -- CP-element group 95: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/$exit
      -- CP-element group 95: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_sources/type_cast_1533/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1527/phi_stmt_1527_req
      -- 
    phi_stmt_1527_req_4358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1527_req_4358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(95), ack => phi_stmt_1527_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(93) & convTransposeA_CP_3548_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1397/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(86) & convTransposeA_CP_3548_elements(89) & convTransposeA_CP_3548_elements(92) & convTransposeA_CP_3548_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1397/merge_stmt_1505_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_1397/merge_stmt_1505_PhiAck/$entry
      -- 
    convTransposeA_CP_3548_elements(97) <= OrReduce(convTransposeA_CP_3548_elements(83) & convTransposeA_CP_3548_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1397/merge_stmt_1505_PhiAck/phi_stmt_1506_ack
      -- 
    phi_stmt_1506_ack_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1506_ack_0, ack => convTransposeA_CP_3548_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1397/merge_stmt_1505_PhiAck/phi_stmt_1513_ack
      -- 
    phi_stmt_1513_ack_4364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1513_ack_0, ack => convTransposeA_CP_3548_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1397/merge_stmt_1505_PhiAck/phi_stmt_1520_ack
      -- 
    phi_stmt_1520_ack_4365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1520_ack_0, ack => convTransposeA_CP_3548_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1397/merge_stmt_1505_PhiAck/phi_stmt_1527_ack
      -- 
    phi_stmt_1527_ack_4366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1527_ack_0, ack => convTransposeA_CP_3548_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1576_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1636_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1612_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/array_obj_ref_1635_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1606_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1572_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1568_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/addr_of_1613_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1617_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/merge_stmt_1505__exit__
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656__entry__
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/ptr_deref_1639_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1397/assign_stmt_1540_to_assign_stmt_1656/type_cast_1644_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1397/merge_stmt_1505_PhiAck/$exit
      -- 
    rr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1576_inst_req_0); -- 
    req_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => array_obj_ref_1612_index_offset_req_1); -- 
    rr_3924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1606_inst_req_0); -- 
    cr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1576_inst_req_1); -- 
    cr_3887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1568_inst_req_1); -- 
    req_4056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => array_obj_ref_1635_index_offset_req_1); -- 
    rr_3896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1572_inst_req_0); -- 
    cr_3901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1572_inst_req_1); -- 
    rr_3882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1568_inst_req_0); -- 
    cr_3929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1606_inst_req_1); -- 
    req_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => addr_of_1636_final_reg_req_1); -- 
    req_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => addr_of_1613_final_reg_req_1); -- 
    cr_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => ptr_deref_1617_load_0_req_1); -- 
    cr_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => ptr_deref_1639_store_0_req_1); -- 
    rr_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1644_inst_req_0); -- 
    cr_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(102), ack => type_cast_1644_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(98) & convTransposeA_CP_3548_elements(99) & convTransposeA_CP_3548_elements(100) & convTransposeA_CP_3548_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  output  delay-element  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	110 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1715/$exit
      -- CP-element group 103: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1721_konst_delay_trans
      -- CP-element group 103: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_req
      -- 
    phi_stmt_1715_req_4401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1715_req_4401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(103), ack => phi_stmt_1715_req_1); -- 
    -- Element group convTransposeA_CP_3548_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => convTransposeA_CP_3548_elements(76), ack => convTransposeA_CP_3548_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Sample/ra
      -- 
    ra_4418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1725_inst_ack_0, ack => convTransposeA_CP_3548_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/Update/ca
      -- 
    ca_4423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1725_inst_ack_1, ack => convTransposeA_CP_3548_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/$exit
      -- CP-element group 106: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/$exit
      -- CP-element group 106: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1725/SplitProtocol/$exit
      -- CP-element group 106: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_req
      -- 
    phi_stmt_1722_req_4424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1722_req_4424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(106), ack => phi_stmt_1722_req_0); -- 
    convTransposeA_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(104) & convTransposeA_CP_3548_elements(105);
      gj_convTransposeA_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Sample/ra
      -- 
    ra_4441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1733_inst_ack_0, ack => convTransposeA_CP_3548_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/Update/ca
      -- 
    ca_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1733_inst_ack_1, ack => convTransposeA_CP_3548_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/$exit
      -- CP-element group 109: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/$exit
      -- CP-element group 109: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1733/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_req
      -- 
    phi_stmt_1728_req_4447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_req_4447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(109), ack => phi_stmt_1728_req_1); -- 
    convTransposeA_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(107) & convTransposeA_CP_3548_elements(108);
      gj_convTransposeA_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1397/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(103) & convTransposeA_CP_3548_elements(106) & convTransposeA_CP_3548_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Sample/ra
      -- 
    ra_4467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_0, ack => convTransposeA_CP_3548_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/Update/ca
      -- 
    ca_4472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_1, ack => convTransposeA_CP_3548_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/$exit
      -- CP-element group 113: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/$exit
      -- CP-element group 113: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_sources/type_cast_1718/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1715/phi_stmt_1715_req
      -- 
    phi_stmt_1715_req_4473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1715_req_4473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(113), ack => phi_stmt_1715_req_0); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(111) & convTransposeA_CP_3548_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Sample/ra
      -- 
    ra_4490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1727_inst_ack_0, ack => convTransposeA_CP_3548_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/Update/ca
      -- 
    ca_4495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1727_inst_ack_1, ack => convTransposeA_CP_3548_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/$exit
      -- CP-element group 116: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/$exit
      -- CP-element group 116: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_sources/type_cast_1727/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1722/phi_stmt_1722_req
      -- 
    phi_stmt_1722_req_4496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1722_req_4496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(116), ack => phi_stmt_1722_req_1); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(114) & convTransposeA_CP_3548_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Sample/ra
      -- 
    ra_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_0, ack => convTransposeA_CP_3548_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/Update/ca
      -- 
    ca_4518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_1, ack => convTransposeA_CP_3548_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/$exit
      -- CP-element group 119: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/$exit
      -- CP-element group 119: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_sources/type_cast_1731/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1728/phi_stmt_1728_req
      -- 
    phi_stmt_1728_req_4519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_req_4519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3548_elements(119), ack => phi_stmt_1728_req_0); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(117) & convTransposeA_CP_3548_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1397/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(113) & convTransposeA_CP_3548_elements(116) & convTransposeA_CP_3548_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1397/merge_stmt_1714_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_1397/merge_stmt_1714_PhiAck/$entry
      -- 
    convTransposeA_CP_3548_elements(121) <= OrReduce(convTransposeA_CP_3548_elements(110) & convTransposeA_CP_3548_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1397/merge_stmt_1714_PhiAck/phi_stmt_1715_ack
      -- 
    phi_stmt_1715_ack_4524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1715_ack_0, ack => convTransposeA_CP_3548_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1397/merge_stmt_1714_PhiAck/phi_stmt_1722_ack
      -- 
    phi_stmt_1722_ack_4525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1722_ack_0, ack => convTransposeA_CP_3548_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1397/merge_stmt_1714_PhiAck/phi_stmt_1728_ack
      -- 
    phi_stmt_1728_ack_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1728_ack_0, ack => convTransposeA_CP_3548_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1397/merge_stmt_1714_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3548_elements(122) & convTransposeA_CP_3548_elements(123) & convTransposeA_CP_3548_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3548_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1634_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1634_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1611_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1611_scaled : std_logic_vector(13 downto 0);
    signal add41_1465 : std_logic_vector(15 downto 0);
    signal add54_1476 : std_logic_vector(15 downto 0);
    signal add73_1587 : std_logic_vector(63 downto 0);
    signal add75_1597 : std_logic_vector(63 downto 0);
    signal add86_1651 : std_logic_vector(31 downto 0);
    signal add93_1669 : std_logic_vector(15 downto 0);
    signal add_1449 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1545 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1612_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1612_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1612_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1612_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1612_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1612_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1635_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1635_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1635_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1635_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1635_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1635_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1614 : std_logic_vector(31 downto 0);
    signal arrayidx82_1637 : std_logic_vector(31 downto 0);
    signal call11_1418 : std_logic_vector(15 downto 0);
    signal call13_1421 : std_logic_vector(15 downto 0);
    signal call14_1424 : std_logic_vector(15 downto 0);
    signal call15_1427 : std_logic_vector(15 downto 0);
    signal call16_1440 : std_logic_vector(15 downto 0);
    signal call18_1452 : std_logic_vector(15 downto 0);
    signal call1_1403 : std_logic_vector(15 downto 0);
    signal call20_1455 : std_logic_vector(15 downto 0);
    signal call22_1458 : std_logic_vector(15 downto 0);
    signal call3_1406 : std_logic_vector(15 downto 0);
    signal call5_1409 : std_logic_vector(15 downto 0);
    signal call7_1412 : std_logic_vector(15 downto 0);
    signal call9_1415 : std_logic_vector(15 downto 0);
    signal call_1400 : std_logic_vector(15 downto 0);
    signal cmp101_1682 : std_logic_vector(0 downto 0);
    signal cmp112_1707 : std_logic_vector(0 downto 0);
    signal cmp_1656 : std_logic_vector(0 downto 0);
    signal conv107_1702 : std_logic_vector(31 downto 0);
    signal conv110_1497 : std_logic_vector(31 downto 0);
    signal conv17_1444 : std_logic_vector(31 downto 0);
    signal conv61_1569 : std_logic_vector(63 downto 0);
    signal conv64_1485 : std_logic_vector(63 downto 0);
    signal conv66_1573 : std_logic_vector(63 downto 0);
    signal conv69_1489 : std_logic_vector(63 downto 0);
    signal conv71_1577 : std_logic_vector(63 downto 0);
    signal conv85_1645 : std_logic_vector(31 downto 0);
    signal conv89_1493 : std_logic_vector(31 downto 0);
    signal conv_1431 : std_logic_vector(31 downto 0);
    signal idxprom81_1630 : std_logic_vector(63 downto 0);
    signal idxprom_1607 : std_logic_vector(63 downto 0);
    signal inc105_1686 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1691 : std_logic_vector(15 downto 0);
    signal inc_1677 : std_logic_vector(15 downto 0);
    signal indvar_1506 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1740 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1728 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1527 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1722 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1520 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1698 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1715 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1513 : std_logic_vector(15 downto 0);
    signal mul50_1560 : std_logic_vector(15 downto 0);
    signal mul72_1582 : std_logic_vector(63 downto 0);
    signal mul74_1592 : std_logic_vector(63 downto 0);
    signal mul_1550 : std_logic_vector(15 downto 0);
    signal ptr_deref_1617_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1617_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1617_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1617_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1617_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1639_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1639_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1437 : std_logic_vector(31 downto 0);
    signal shr111126_1503 : std_logic_vector(31 downto 0);
    signal shr80_1624 : std_logic_vector(63 downto 0);
    signal shr_1603 : std_logic_vector(31 downto 0);
    signal sub44_1555 : std_logic_vector(15 downto 0);
    signal sub57_1481 : std_logic_vector(15 downto 0);
    signal sub58_1565 : std_logic_vector(15 downto 0);
    signal sub_1470 : std_logic_vector(15 downto 0);
    signal tmp1_1540 : std_logic_vector(31 downto 0);
    signal tmp78_1618 : std_logic_vector(63 downto 0);
    signal type_cast_1435_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1463_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1474_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1501_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1512_wire : std_logic_vector(31 downto 0);
    signal type_cast_1517_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1519_wire : std_logic_vector(15 downto 0);
    signal type_cast_1524_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1526_wire : std_logic_vector(15 downto 0);
    signal type_cast_1531_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1533_wire : std_logic_vector(15 downto 0);
    signal type_cast_1538_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1601_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1622_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1628_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1667_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1675_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1695_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1718_wire : std_logic_vector(15 downto 0);
    signal type_cast_1721_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1725_wire : std_logic_vector(15 downto 0);
    signal type_cast_1727_wire : std_logic_vector(15 downto 0);
    signal type_cast_1731_wire : std_logic_vector(15 downto 0);
    signal type_cast_1733_wire : std_logic_vector(15 downto 0);
    signal type_cast_1738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1746_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1612_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1612_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1612_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1612_resized_base_address <= "00000000000000";
    array_obj_ref_1635_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1635_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1635_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1635_resized_base_address <= "00000000000000";
    ptr_deref_1617_word_offset_0 <= "00000000000000";
    ptr_deref_1639_word_offset_0 <= "00000000000000";
    type_cast_1435_wire_constant <= "00000000000000000000000000010000";
    type_cast_1463_wire_constant <= "1111111111111111";
    type_cast_1474_wire_constant <= "1111111111111111";
    type_cast_1501_wire_constant <= "00000000000000000000000000000010";
    type_cast_1510_wire_constant <= "00000000000000000000000000000000";
    type_cast_1517_wire_constant <= "0000000000000000";
    type_cast_1524_wire_constant <= "0000000000000000";
    type_cast_1531_wire_constant <= "0000000000000000";
    type_cast_1538_wire_constant <= "00000000000000000000000000000100";
    type_cast_1601_wire_constant <= "00000000000000000000000000000010";
    type_cast_1622_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1628_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1649_wire_constant <= "00000000000000000000000000000100";
    type_cast_1667_wire_constant <= "0000000000000100";
    type_cast_1675_wire_constant <= "0000000000000001";
    type_cast_1695_wire_constant <= "0000000000000000";
    type_cast_1721_wire_constant <= "0000000000000000";
    type_cast_1738_wire_constant <= "00000000000000000000000000000001";
    type_cast_1746_wire_constant <= "0000000000000001";
    phi_stmt_1506: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1510_wire_constant & type_cast_1512_wire;
      req <= phi_stmt_1506_req_0 & phi_stmt_1506_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1506",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1506_ack_0,
          idata => idata,
          odata => indvar_1506,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1506
    phi_stmt_1513: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1517_wire_constant & type_cast_1519_wire;
      req <= phi_stmt_1513_req_0 & phi_stmt_1513_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1513",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1513_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1513,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1513
    phi_stmt_1520: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1524_wire_constant & type_cast_1526_wire;
      req <= phi_stmt_1520_req_0 & phi_stmt_1520_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1520",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1520_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1520,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1520
    phi_stmt_1527: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1531_wire_constant & type_cast_1533_wire;
      req <= phi_stmt_1527_req_0 & phi_stmt_1527_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1527",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1527_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1527,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1527
    phi_stmt_1715: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1718_wire & type_cast_1721_wire_constant;
      req <= phi_stmt_1715_req_0 & phi_stmt_1715_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1715",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1715_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1715,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1715
    phi_stmt_1722: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1725_wire & type_cast_1727_wire;
      req <= phi_stmt_1722_req_0 & phi_stmt_1722_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1722",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1722_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1722,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1722
    phi_stmt_1728: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1731_wire & type_cast_1733_wire;
      req <= phi_stmt_1728_req_0 & phi_stmt_1728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1728",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1728_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1728
    -- flow-through select operator MUX_1697_inst
    input_dim1x_x2_1698 <= type_cast_1695_wire_constant when (cmp101_1682(0) /=  '0') else inc_1677;
    addr_of_1613_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1613_final_reg_req_0;
      addr_of_1613_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1613_final_reg_req_1;
      addr_of_1613_final_reg_ack_1<= rack(0);
      addr_of_1613_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1613_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1612_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1636_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1636_final_reg_req_0;
      addr_of_1636_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1636_final_reg_req_1;
      addr_of_1636_final_reg_ack_1<= rack(0);
      addr_of_1636_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1636_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1635_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1430_inst_req_0;
      type_cast_1430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1430_inst_req_1;
      type_cast_1430_inst_ack_1<= rack(0);
      type_cast_1430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1443_inst_req_0;
      type_cast_1443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1443_inst_req_1;
      type_cast_1443_inst_ack_1<= rack(0);
      type_cast_1443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1484_inst_req_0;
      type_cast_1484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1484_inst_req_1;
      type_cast_1484_inst_ack_1<= rack(0);
      type_cast_1484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1488_inst_req_0;
      type_cast_1488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1488_inst_req_1;
      type_cast_1488_inst_ack_1<= rack(0);
      type_cast_1488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1492_inst_req_0;
      type_cast_1492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1492_inst_req_1;
      type_cast_1492_inst_ack_1<= rack(0);
      type_cast_1492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1496_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1496_inst_req_0;
      type_cast_1496_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1496_inst_req_1;
      type_cast_1496_inst_ack_1<= rack(0);
      type_cast_1496_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1496_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1400,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1497,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1512_inst_req_0;
      type_cast_1512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1512_inst_req_1;
      type_cast_1512_inst_ack_1<= rack(0);
      type_cast_1512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1512_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1519_inst_req_0;
      type_cast_1519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1519_inst_req_1;
      type_cast_1519_inst_ack_1<= rack(0);
      type_cast_1519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1519_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1526_inst_req_0;
      type_cast_1526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1526_inst_req_1;
      type_cast_1526_inst_ack_1<= rack(0);
      type_cast_1526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1526_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1722,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1526_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1533_inst_req_0;
      type_cast_1533_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1533_inst_req_1;
      type_cast_1533_inst_ack_1<= rack(0);
      type_cast_1533_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1533_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1533_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1568_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1568_inst_req_0;
      type_cast_1568_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1568_inst_req_1;
      type_cast_1568_inst_ack_1<= rack(0);
      type_cast_1568_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1568_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1513,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1569,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1572_inst_req_0;
      type_cast_1572_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1572_inst_req_1;
      type_cast_1572_inst_ack_1<= rack(0);
      type_cast_1572_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1572_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1573,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1576_inst_req_0;
      type_cast_1576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1576_inst_req_1;
      type_cast_1576_inst_ack_1<= rack(0);
      type_cast_1576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1606_inst_req_0;
      type_cast_1606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1606_inst_req_1;
      type_cast_1606_inst_ack_1<= rack(0);
      type_cast_1606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1644_inst_req_0;
      type_cast_1644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1644_inst_req_1;
      type_cast_1644_inst_ack_1<= rack(0);
      type_cast_1644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1513,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1685_inst_req_0;
      type_cast_1685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1685_inst_req_1;
      type_cast_1685_inst_ack_1<= rack(0);
      type_cast_1685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1682,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1701_inst_req_0;
      type_cast_1701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1701_inst_req_1;
      type_cast_1701_inst_ack_1<= rack(0);
      type_cast_1701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1718_inst_req_0;
      type_cast_1718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1718_inst_req_1;
      type_cast_1718_inst_ack_1<= rack(0);
      type_cast_1718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1718_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1725_inst_req_0;
      type_cast_1725_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1725_inst_req_1;
      type_cast_1725_inst_ack_1<= rack(0);
      type_cast_1725_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1725_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1725_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1727_inst_req_0;
      type_cast_1727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1727_inst_req_1;
      type_cast_1727_inst_ack_1<= rack(0);
      type_cast_1727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1727_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1731_inst_req_0;
      type_cast_1731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1731_inst_req_1;
      type_cast_1731_inst_ack_1<= rack(0);
      type_cast_1731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1527,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1731_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1733_inst_req_0;
      type_cast_1733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1733_inst_req_1;
      type_cast_1733_inst_ack_1<= rack(0);
      type_cast_1733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1733_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1612_index_1_rename
    process(R_idxprom_1611_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1611_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1611_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1612_index_1_resize
    process(idxprom_1607) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1607;
      ov := iv(13 downto 0);
      R_idxprom_1611_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1612_root_address_inst
    process(array_obj_ref_1612_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1612_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1612_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1635_index_1_rename
    process(R_idxprom81_1634_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1634_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1634_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1635_index_1_resize
    process(idxprom81_1630) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1630;
      ov := iv(13 downto 0);
      R_idxprom81_1634_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1635_root_address_inst
    process(array_obj_ref_1635_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1635_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1635_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1617_addr_0
    process(ptr_deref_1617_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1617_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1617_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1617_base_resize
    process(arrayidx77_1614) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1614;
      ov := iv(13 downto 0);
      ptr_deref_1617_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1617_gather_scatter
    process(ptr_deref_1617_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1617_data_0;
      ov(63 downto 0) := iv;
      tmp78_1618 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1617_root_address_inst
    process(ptr_deref_1617_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1617_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1617_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_addr_0
    process(ptr_deref_1639_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1639_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1639_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_base_resize
    process(arrayidx82_1637) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1637;
      ov := iv(13 downto 0);
      ptr_deref_1639_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_gather_scatter
    process(tmp78_1618) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1618;
      ov(63 downto 0) := iv;
      ptr_deref_1639_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_root_address_inst
    process(ptr_deref_1639_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1639_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1639_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1657_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1656;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1657_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1657_branch_req_0,
          ack0 => if_stmt_1657_branch_ack_0,
          ack1 => if_stmt_1657_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1708_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1707;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1708_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1708_branch_req_0,
          ack0 => if_stmt_1708_branch_ack_0,
          ack1 => if_stmt_1708_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1464_inst
    process(call7_1412) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1412, type_cast_1463_wire_constant, tmp_var);
      add41_1465 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1475_inst
    process(call9_1415) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1415, type_cast_1474_wire_constant, tmp_var);
      add54_1476 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1554_inst
    process(sub_1470, mul_1550) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1470, mul_1550, tmp_var);
      sub44_1555 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1564_inst
    process(sub57_1481, mul50_1560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1481, mul50_1560, tmp_var);
      sub58_1565 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1668_inst
    process(input_dim2x_x1_1513) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1513, type_cast_1667_wire_constant, tmp_var);
      add93_1669 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1676_inst
    process(input_dim1x_x1_1520) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1520, type_cast_1675_wire_constant, tmp_var);
      inc_1677 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1690_inst
    process(inc105_1686, input_dim0x_x2_1527) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1686, input_dim0x_x2_1527, tmp_var);
      inc105x_xinput_dim0x_x2_1691 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1544_inst
    process(add_1449, tmp1_1540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1449, tmp1_1540, tmp_var);
      add_src_0x_x0_1545 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1650_inst
    process(conv85_1645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1645, type_cast_1649_wire_constant, tmp_var);
      add86_1651 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1739_inst
    process(indvar_1506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1506, type_cast_1738_wire_constant, tmp_var);
      indvarx_xnext_1740 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1586_inst
    process(mul72_1582, conv66_1573) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1582, conv66_1573, tmp_var);
      add73_1587 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1596_inst
    process(mul74_1592, conv61_1569) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1592, conv61_1569, tmp_var);
      add75_1597 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1629_inst
    process(shr80_1624) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1624, type_cast_1628_wire_constant, tmp_var);
      idxprom81_1630 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1681_inst
    process(inc_1677, call1_1403) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1677, call1_1403, tmp_var);
      cmp101_1682 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1706_inst
    process(conv107_1702, shr111126_1503) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1702, shr111126_1503, tmp_var);
      cmp112_1707 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1502_inst
    process(conv110_1497) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1497, type_cast_1501_wire_constant, tmp_var);
      shr111126_1503 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1602_inst
    process(add_src_0x_x0_1545) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1545, type_cast_1601_wire_constant, tmp_var);
      shr_1603 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1623_inst
    process(add75_1597) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1597, type_cast_1622_wire_constant, tmp_var);
      shr80_1624 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1549_inst
    process(input_dim0x_x2_1527, call13_1421) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1527, call13_1421, tmp_var);
      mul_1550 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1559_inst
    process(input_dim1x_x1_1520, call13_1421) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1520, call13_1421, tmp_var);
      mul50_1560 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1539_inst
    process(indvar_1506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1506, type_cast_1538_wire_constant, tmp_var);
      tmp1_1540 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1581_inst
    process(conv71_1577, conv69_1489) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1577, conv69_1489, tmp_var);
      mul72_1582 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1591_inst
    process(add73_1587, conv64_1485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1587, conv64_1485, tmp_var);
      mul74_1592 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1448_inst
    process(shl_1437, conv17_1444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1437, conv17_1444, tmp_var);
      add_1449 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1436_inst
    process(conv_1431) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1431, type_cast_1435_wire_constant, tmp_var);
      shl_1437 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1469_inst
    process(add41_1465, call14_1424) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1465, call14_1424, tmp_var);
      sub_1470 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1480_inst
    process(add54_1476, call14_1424) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1476, call14_1424, tmp_var);
      sub57_1481 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1655_inst
    process(add86_1651, conv89_1493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1651, conv89_1493, tmp_var);
      cmp_1656 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1612_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1611_scaled;
      array_obj_ref_1612_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1612_index_offset_req_0;
      array_obj_ref_1612_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1612_index_offset_req_1;
      array_obj_ref_1612_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1635_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1634_scaled;
      array_obj_ref_1635_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1635_index_offset_req_0;
      array_obj_ref_1635_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1635_index_offset_req_1;
      array_obj_ref_1635_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1617_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1617_load_0_req_0;
      ptr_deref_1617_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1617_load_0_req_1;
      ptr_deref_1617_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1617_word_address_0;
      ptr_deref_1617_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1639_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1639_store_0_req_0;
      ptr_deref_1639_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1639_store_0_req_1;
      ptr_deref_1639_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1639_word_address_0;
      data_in <= ptr_deref_1639_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1420_inst RPIPE_Block0_start_1423_inst RPIPE_Block0_start_1426_inst RPIPE_Block0_start_1457_inst RPIPE_Block0_start_1439_inst RPIPE_Block0_start_1451_inst RPIPE_Block0_start_1454_inst RPIPE_Block0_start_1417_inst RPIPE_Block0_start_1414_inst RPIPE_Block0_start_1411_inst RPIPE_Block0_start_1408_inst RPIPE_Block0_start_1405_inst RPIPE_Block0_start_1402_inst RPIPE_Block0_start_1399_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1420_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1423_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1426_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1457_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1439_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1451_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1454_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1417_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1414_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1411_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1408_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1405_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1402_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1399_inst_req_0;
      RPIPE_Block0_start_1420_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1423_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1426_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1457_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1439_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1451_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1454_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1417_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1414_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1411_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1408_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1405_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1402_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1399_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1420_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1423_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1426_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1457_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1439_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1451_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1454_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1417_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1414_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1411_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1408_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1405_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1402_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1399_inst_req_1;
      RPIPE_Block0_start_1420_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1423_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1426_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1457_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1439_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1451_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1454_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1417_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1414_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1411_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1408_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1405_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1402_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1399_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call13_1421 <= data_out(223 downto 208);
      call14_1424 <= data_out(207 downto 192);
      call15_1427 <= data_out(191 downto 176);
      call22_1458 <= data_out(175 downto 160);
      call16_1440 <= data_out(159 downto 144);
      call18_1452 <= data_out(143 downto 128);
      call20_1455 <= data_out(127 downto 112);
      call11_1418 <= data_out(111 downto 96);
      call9_1415 <= data_out(95 downto 80);
      call7_1412 <= data_out(79 downto 64);
      call5_1409 <= data_out(63 downto 48);
      call3_1406 <= data_out(47 downto 32);
      call1_1403 <= data_out(31 downto 16);
      call_1400 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1744_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1744_inst_req_0;
      WPIPE_Block0_done_1744_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1744_inst_req_1;
      WPIPE_Block0_done_1744_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1746_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4543_start: Boolean;
  signal convTransposeB_CP_4543_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2005_inst_req_0 : boolean;
  signal addr_of_1997_final_reg_req_0 : boolean;
  signal ptr_deref_2000_store_0_req_0 : boolean;
  signal array_obj_ref_1996_index_offset_ack_0 : boolean;
  signal array_obj_ref_1996_index_offset_ack_1 : boolean;
  signal addr_of_1997_final_reg_ack_0 : boolean;
  signal type_cast_2005_inst_ack_0 : boolean;
  signal if_stmt_2018_branch_ack_1 : boolean;
  signal if_stmt_2018_branch_req_0 : boolean;
  signal ptr_deref_2000_store_0_req_1 : boolean;
  signal type_cast_2005_inst_ack_1 : boolean;
  signal ptr_deref_2000_store_0_ack_1 : boolean;
  signal array_obj_ref_1996_index_offset_req_1 : boolean;
  signal ptr_deref_2000_store_0_ack_0 : boolean;
  signal addr_of_1997_final_reg_req_1 : boolean;
  signal addr_of_1997_final_reg_ack_1 : boolean;
  signal array_obj_ref_1996_index_offset_req_0 : boolean;
  signal RPIPE_Block1_start_1755_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1755_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1755_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1755_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1758_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1758_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1758_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1758_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1761_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1761_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1761_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1761_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1764_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1764_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1764_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1764_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1767_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1767_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1767_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1767_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1770_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1770_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1770_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1770_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1773_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1773_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1773_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1773_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1776_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1776_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1776_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1776_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1779_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1779_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1779_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1779_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1782_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1782_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1782_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1782_inst_ack_1 : boolean;
  signal type_cast_1786_inst_req_0 : boolean;
  signal type_cast_1786_inst_ack_0 : boolean;
  signal type_cast_1786_inst_req_1 : boolean;
  signal type_cast_1786_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1795_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1795_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1795_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1795_inst_ack_1 : boolean;
  signal type_cast_1799_inst_req_0 : boolean;
  signal type_cast_1799_inst_ack_0 : boolean;
  signal type_cast_1799_inst_req_1 : boolean;
  signal type_cast_1799_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1807_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1807_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1807_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1807_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1810_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1810_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1810_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1810_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1813_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1813_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1813_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1813_inst_ack_1 : boolean;
  signal type_cast_1846_inst_req_0 : boolean;
  signal type_cast_1846_inst_ack_0 : boolean;
  signal type_cast_1846_inst_req_1 : boolean;
  signal type_cast_1846_inst_ack_1 : boolean;
  signal type_cast_1850_inst_req_0 : boolean;
  signal type_cast_1850_inst_ack_0 : boolean;
  signal type_cast_1850_inst_req_1 : boolean;
  signal type_cast_1850_inst_ack_1 : boolean;
  signal type_cast_1854_inst_req_0 : boolean;
  signal type_cast_1854_inst_ack_0 : boolean;
  signal type_cast_1854_inst_req_1 : boolean;
  signal type_cast_1854_inst_ack_1 : boolean;
  signal type_cast_1858_inst_req_0 : boolean;
  signal type_cast_1858_inst_ack_0 : boolean;
  signal type_cast_1858_inst_req_1 : boolean;
  signal type_cast_1858_inst_ack_1 : boolean;
  signal type_cast_1929_inst_req_0 : boolean;
  signal type_cast_1929_inst_ack_0 : boolean;
  signal type_cast_1929_inst_req_1 : boolean;
  signal type_cast_1929_inst_ack_1 : boolean;
  signal type_cast_1933_inst_req_0 : boolean;
  signal type_cast_1933_inst_ack_0 : boolean;
  signal type_cast_1933_inst_req_1 : boolean;
  signal type_cast_1933_inst_ack_1 : boolean;
  signal type_cast_1937_inst_req_0 : boolean;
  signal type_cast_1937_inst_ack_0 : boolean;
  signal type_cast_1937_inst_req_1 : boolean;
  signal type_cast_1937_inst_ack_1 : boolean;
  signal type_cast_1967_inst_req_0 : boolean;
  signal type_cast_1967_inst_ack_0 : boolean;
  signal type_cast_1967_inst_req_1 : boolean;
  signal type_cast_1967_inst_ack_1 : boolean;
  signal type_cast_2005_inst_req_1 : boolean;
  signal array_obj_ref_1973_index_offset_req_0 : boolean;
  signal array_obj_ref_1973_index_offset_ack_0 : boolean;
  signal array_obj_ref_1973_index_offset_req_1 : boolean;
  signal array_obj_ref_1973_index_offset_ack_1 : boolean;
  signal addr_of_1974_final_reg_req_0 : boolean;
  signal addr_of_1974_final_reg_ack_0 : boolean;
  signal addr_of_1974_final_reg_req_1 : boolean;
  signal addr_of_1974_final_reg_ack_1 : boolean;
  signal ptr_deref_1978_load_0_req_0 : boolean;
  signal ptr_deref_1978_load_0_ack_0 : boolean;
  signal ptr_deref_1978_load_0_req_1 : boolean;
  signal ptr_deref_1978_load_0_ack_1 : boolean;
  signal if_stmt_2018_branch_ack_0 : boolean;
  signal type_cast_2046_inst_req_0 : boolean;
  signal type_cast_2046_inst_ack_0 : boolean;
  signal type_cast_2046_inst_req_1 : boolean;
  signal type_cast_2046_inst_ack_1 : boolean;
  signal type_cast_2062_inst_req_0 : boolean;
  signal type_cast_2062_inst_ack_0 : boolean;
  signal type_cast_2062_inst_req_1 : boolean;
  signal type_cast_2062_inst_ack_1 : boolean;
  signal if_stmt_2069_branch_req_0 : boolean;
  signal if_stmt_2069_branch_ack_1 : boolean;
  signal if_stmt_2069_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2105_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2105_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2105_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2105_inst_ack_1 : boolean;
  signal type_cast_1892_inst_req_0 : boolean;
  signal type_cast_1892_inst_ack_0 : boolean;
  signal type_cast_1892_inst_req_1 : boolean;
  signal type_cast_1892_inst_ack_1 : boolean;
  signal phi_stmt_1889_req_0 : boolean;
  signal phi_stmt_1882_req_0 : boolean;
  signal phi_stmt_1875_req_0 : boolean;
  signal phi_stmt_1868_req_0 : boolean;
  signal type_cast_1894_inst_req_0 : boolean;
  signal type_cast_1894_inst_ack_0 : boolean;
  signal type_cast_1894_inst_req_1 : boolean;
  signal type_cast_1894_inst_ack_1 : boolean;
  signal phi_stmt_1889_req_1 : boolean;
  signal type_cast_1888_inst_req_0 : boolean;
  signal type_cast_1888_inst_ack_0 : boolean;
  signal type_cast_1888_inst_req_1 : boolean;
  signal type_cast_1888_inst_ack_1 : boolean;
  signal phi_stmt_1882_req_1 : boolean;
  signal type_cast_1881_inst_req_0 : boolean;
  signal type_cast_1881_inst_ack_0 : boolean;
  signal type_cast_1881_inst_req_1 : boolean;
  signal type_cast_1881_inst_ack_1 : boolean;
  signal phi_stmt_1875_req_1 : boolean;
  signal type_cast_1874_inst_req_0 : boolean;
  signal type_cast_1874_inst_ack_0 : boolean;
  signal type_cast_1874_inst_req_1 : boolean;
  signal type_cast_1874_inst_ack_1 : boolean;
  signal phi_stmt_1868_req_1 : boolean;
  signal phi_stmt_1868_ack_0 : boolean;
  signal phi_stmt_1875_ack_0 : boolean;
  signal phi_stmt_1882_ack_0 : boolean;
  signal phi_stmt_1889_ack_0 : boolean;
  signal type_cast_2094_inst_req_0 : boolean;
  signal type_cast_2094_inst_ack_0 : boolean;
  signal type_cast_2094_inst_req_1 : boolean;
  signal type_cast_2094_inst_ack_1 : boolean;
  signal phi_stmt_2089_req_1 : boolean;
  signal type_cast_2086_inst_req_0 : boolean;
  signal type_cast_2086_inst_ack_0 : boolean;
  signal type_cast_2086_inst_req_1 : boolean;
  signal type_cast_2086_inst_ack_1 : boolean;
  signal phi_stmt_2083_req_0 : boolean;
  signal phi_stmt_2076_req_1 : boolean;
  signal type_cast_2092_inst_req_0 : boolean;
  signal type_cast_2092_inst_ack_0 : boolean;
  signal type_cast_2092_inst_req_1 : boolean;
  signal type_cast_2092_inst_ack_1 : boolean;
  signal phi_stmt_2089_req_0 : boolean;
  signal type_cast_2088_inst_req_0 : boolean;
  signal type_cast_2088_inst_ack_0 : boolean;
  signal type_cast_2088_inst_req_1 : boolean;
  signal type_cast_2088_inst_ack_1 : boolean;
  signal phi_stmt_2083_req_1 : boolean;
  signal type_cast_2079_inst_req_0 : boolean;
  signal type_cast_2079_inst_ack_0 : boolean;
  signal type_cast_2079_inst_req_1 : boolean;
  signal type_cast_2079_inst_ack_1 : boolean;
  signal phi_stmt_2076_req_0 : boolean;
  signal phi_stmt_2076_ack_0 : boolean;
  signal phi_stmt_2083_ack_0 : boolean;
  signal phi_stmt_2089_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4543_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4543_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4543_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4543_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4543: Block -- control-path 
    signal convTransposeB_CP_4543_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4543_elements(0) <= convTransposeB_CP_4543_start;
    convTransposeB_CP_4543_symbol <= convTransposeB_CP_4543_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1753/$entry
      -- CP-element group 0: 	 branch_block_stmt_1753/branch_block_stmt_1753__entry__
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814__entry__
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/$entry
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Update/cr
      -- 
    rr_4591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(0), ack => RPIPE_Block1_start_1755_inst_req_0); -- 
    cr_4736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(0), ack => type_cast_1786_inst_req_1); -- 
    cr_4764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(0), ack => type_cast_1799_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1753/merge_stmt_2075__exit__
      -- CP-element group 1: 	 branch_block_stmt_1753/assign_stmt_2101__entry__
      -- CP-element group 1: 	 branch_block_stmt_1753/assign_stmt_2101__exit__
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1753/assign_stmt_2101/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/assign_stmt_2101/$exit
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/cr
      -- 
    rr_5292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1894_inst_req_0); -- 
    cr_5297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1894_inst_req_1); -- 
    rr_5315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1888_inst_req_0); -- 
    cr_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1888_inst_req_1); -- 
    rr_5338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1881_inst_req_0); -- 
    cr_5343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1881_inst_req_1); -- 
    rr_5361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1874_inst_req_0); -- 
    cr_5366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(1), ack => type_cast_1874_inst_req_1); -- 
    convTransposeB_CP_4543_elements(1) <= convTransposeB_CP_4543_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Update/cr
      -- 
    ra_4592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1755_inst_ack_0, ack => convTransposeB_CP_4543_elements(2)); -- 
    cr_4596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(2), ack => RPIPE_Block1_start_1755_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1755_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Sample/rr
      -- 
    ca_4597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1755_inst_ack_1, ack => convTransposeB_CP_4543_elements(3)); -- 
    rr_4605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(3), ack => RPIPE_Block1_start_1758_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Update/cr
      -- 
    ra_4606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1758_inst_ack_0, ack => convTransposeB_CP_4543_elements(4)); -- 
    cr_4610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(4), ack => RPIPE_Block1_start_1758_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1758_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Sample/rr
      -- 
    ca_4611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1758_inst_ack_1, ack => convTransposeB_CP_4543_elements(5)); -- 
    rr_4619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(5), ack => RPIPE_Block1_start_1761_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Update/cr
      -- 
    ra_4620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1761_inst_ack_0, ack => convTransposeB_CP_4543_elements(6)); -- 
    cr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(6), ack => RPIPE_Block1_start_1761_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1761_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Sample/rr
      -- 
    ca_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1761_inst_ack_1, ack => convTransposeB_CP_4543_elements(7)); -- 
    rr_4633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(7), ack => RPIPE_Block1_start_1764_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Update/cr
      -- 
    ra_4634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1764_inst_ack_0, ack => convTransposeB_CP_4543_elements(8)); -- 
    cr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(8), ack => RPIPE_Block1_start_1764_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1764_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Sample/rr
      -- 
    ca_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1764_inst_ack_1, ack => convTransposeB_CP_4543_elements(9)); -- 
    rr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(9), ack => RPIPE_Block1_start_1767_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Update/cr
      -- 
    ra_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1767_inst_ack_0, ack => convTransposeB_CP_4543_elements(10)); -- 
    cr_4652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(10), ack => RPIPE_Block1_start_1767_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1767_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Sample/rr
      -- 
    ca_4653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1767_inst_ack_1, ack => convTransposeB_CP_4543_elements(11)); -- 
    rr_4661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(11), ack => RPIPE_Block1_start_1770_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Update/cr
      -- 
    ra_4662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1770_inst_ack_0, ack => convTransposeB_CP_4543_elements(12)); -- 
    cr_4666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(12), ack => RPIPE_Block1_start_1770_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1770_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Sample/rr
      -- 
    ca_4667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1770_inst_ack_1, ack => convTransposeB_CP_4543_elements(13)); -- 
    rr_4675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(13), ack => RPIPE_Block1_start_1773_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Update/cr
      -- 
    ra_4676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1773_inst_ack_0, ack => convTransposeB_CP_4543_elements(14)); -- 
    cr_4680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(14), ack => RPIPE_Block1_start_1773_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1773_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Sample/rr
      -- 
    ca_4681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1773_inst_ack_1, ack => convTransposeB_CP_4543_elements(15)); -- 
    rr_4689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(15), ack => RPIPE_Block1_start_1776_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Update/cr
      -- 
    ra_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1776_inst_ack_0, ack => convTransposeB_CP_4543_elements(16)); -- 
    cr_4694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(16), ack => RPIPE_Block1_start_1776_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1776_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Sample/rr
      -- 
    ca_4695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1776_inst_ack_1, ack => convTransposeB_CP_4543_elements(17)); -- 
    rr_4703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(17), ack => RPIPE_Block1_start_1779_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Update/cr
      -- 
    ra_4704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1779_inst_ack_0, ack => convTransposeB_CP_4543_elements(18)); -- 
    cr_4708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(18), ack => RPIPE_Block1_start_1779_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1779_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Sample/rr
      -- 
    ca_4709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1779_inst_ack_1, ack => convTransposeB_CP_4543_elements(19)); -- 
    rr_4717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(19), ack => RPIPE_Block1_start_1782_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Update/cr
      -- 
    ra_4718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1782_inst_ack_0, ack => convTransposeB_CP_4543_elements(20)); -- 
    cr_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(20), ack => RPIPE_Block1_start_1782_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1782_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Sample/rr
      -- 
    ca_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1782_inst_ack_1, ack => convTransposeB_CP_4543_elements(21)); -- 
    rr_4731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(21), ack => type_cast_1786_inst_req_0); -- 
    rr_4745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(21), ack => RPIPE_Block1_start_1795_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Sample/ra
      -- 
    ra_4732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1786_inst_ack_0, ack => convTransposeB_CP_4543_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1786_Update/ca
      -- 
    ca_4737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1786_inst_ack_1, ack => convTransposeB_CP_4543_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Update/cr
      -- 
    ra_4746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1795_inst_ack_0, ack => convTransposeB_CP_4543_elements(24)); -- 
    cr_4750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(24), ack => RPIPE_Block1_start_1795_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1795_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Sample/rr
      -- 
    ca_4751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1795_inst_ack_1, ack => convTransposeB_CP_4543_elements(25)); -- 
    rr_4759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(25), ack => type_cast_1799_inst_req_0); -- 
    rr_4773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(25), ack => RPIPE_Block1_start_1807_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Sample/ra
      -- 
    ra_4760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_0, ack => convTransposeB_CP_4543_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/type_cast_1799_Update/ca
      -- 
    ca_4765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_1, ack => convTransposeB_CP_4543_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Update/cr
      -- 
    ra_4774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1807_inst_ack_0, ack => convTransposeB_CP_4543_elements(28)); -- 
    cr_4778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(28), ack => RPIPE_Block1_start_1807_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1807_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Sample/rr
      -- 
    ca_4779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1807_inst_ack_1, ack => convTransposeB_CP_4543_elements(29)); -- 
    rr_4787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(29), ack => RPIPE_Block1_start_1810_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Update/cr
      -- 
    ra_4788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1810_inst_ack_0, ack => convTransposeB_CP_4543_elements(30)); -- 
    cr_4792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(30), ack => RPIPE_Block1_start_1810_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1810_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Sample/rr
      -- 
    ca_4793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1810_inst_ack_1, ack => convTransposeB_CP_4543_elements(31)); -- 
    rr_4801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(31), ack => RPIPE_Block1_start_1813_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Update/cr
      -- 
    ra_4802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1813_inst_ack_0, ack => convTransposeB_CP_4543_elements(32)); -- 
    cr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(32), ack => RPIPE_Block1_start_1813_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/RPIPE_Block1_start_1813_Update/ca
      -- 
    ca_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1813_inst_ack_1, ack => convTransposeB_CP_4543_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814__exit__
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865__entry__
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1756_to_assign_stmt_1814/$exit
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Update/cr
      -- 
    rr_4818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1846_inst_req_0); -- 
    cr_4823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1846_inst_req_1); -- 
    rr_4832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1850_inst_req_0); -- 
    cr_4837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1850_inst_req_1); -- 
    rr_4846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1854_inst_req_0); -- 
    cr_4851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1854_inst_req_1); -- 
    rr_4860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1858_inst_req_0); -- 
    cr_4865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(34), ack => type_cast_1858_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(23) & convTransposeB_CP_4543_elements(27) & convTransposeB_CP_4543_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Sample/ra
      -- 
    ra_4819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1846_inst_ack_0, ack => convTransposeB_CP_4543_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1846_Update/ca
      -- 
    ca_4824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1846_inst_ack_1, ack => convTransposeB_CP_4543_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Sample/ra
      -- 
    ra_4833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_0, ack => convTransposeB_CP_4543_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1850_Update/ca
      -- 
    ca_4838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_1, ack => convTransposeB_CP_4543_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Sample/ra
      -- 
    ra_4847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1854_inst_ack_0, ack => convTransposeB_CP_4543_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1854_Update/ca
      -- 
    ca_4852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1854_inst_ack_1, ack => convTransposeB_CP_4543_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Sample/ra
      -- 
    ra_4861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_0, ack => convTransposeB_CP_4543_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/type_cast_1858_Update/ca
      -- 
    ca_4866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_1, ack => convTransposeB_CP_4543_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865__exit__
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1753/assign_stmt_1821_to_assign_stmt_1865/$exit
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1882/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1875/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1868/$entry
      -- CP-element group 43: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$entry
      -- 
    rr_5242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(43), ack => type_cast_1892_inst_req_0); -- 
    cr_5247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(43), ack => type_cast_1892_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(36) & convTransposeB_CP_4543_elements(38) & convTransposeB_CP_4543_elements(40) & convTransposeB_CP_4543_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Sample/ra
      -- 
    ra_4878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1929_inst_ack_0, ack => convTransposeB_CP_4543_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Update/ca
      -- 
    ca_4883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1929_inst_ack_1, ack => convTransposeB_CP_4543_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Sample/ra
      -- 
    ra_4892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_0, ack => convTransposeB_CP_4543_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Update/ca
      -- 
    ca_4897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_1, ack => convTransposeB_CP_4543_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Sample/ra
      -- 
    ra_4906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_0, ack => convTransposeB_CP_4543_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Update/ca
      -- 
    ca_4911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_1, ack => convTransposeB_CP_4543_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Sample/ra
      -- 
    ra_4920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1967_inst_ack_0, ack => convTransposeB_CP_4543_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Sample/req
      -- 
    ca_4925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1967_inst_ack_1, ack => convTransposeB_CP_4543_elements(51)); -- 
    req_4950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(51), ack => array_obj_ref_1973_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Sample/ack
      -- 
    ack_4951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1973_index_offset_ack_0, ack => convTransposeB_CP_4543_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_request/req
      -- 
    ack_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1973_index_offset_ack_1, ack => convTransposeB_CP_4543_elements(53)); -- 
    req_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(53), ack => addr_of_1974_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_request/ack
      -- 
    ack_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1974_final_reg_ack_0, ack => convTransposeB_CP_4543_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/word_access_start/word_0/rr
      -- 
    ack_4971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1974_final_reg_ack_1, ack => convTransposeB_CP_4543_elements(55)); -- 
    rr_5004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(55), ack => ptr_deref_1978_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Sample/word_access_start/word_0/ra
      -- 
    ra_5005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1978_load_0_ack_0, ack => convTransposeB_CP_4543_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/ptr_deref_1978_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/ptr_deref_1978_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/ptr_deref_1978_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/ptr_deref_1978_Merge/merge_ack
      -- 
    ca_5016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1978_load_0_ack_1, ack => convTransposeB_CP_4543_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_index_resize_1/index_resize_ack
      -- 
    req_5046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(58), ack => array_obj_ref_1996_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(45) & convTransposeB_CP_4543_elements(47) & convTransposeB_CP_4543_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Sample/$exit
      -- 
    ack_5047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1996_index_offset_ack_0, ack => convTransposeB_CP_4543_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_request/req
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_offset_calculated
      -- 
    ack_5052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1996_index_offset_ack_1, ack => convTransposeB_CP_4543_elements(60)); -- 
    req_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(60), ack => addr_of_1997_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_request/ack
      -- CP-element group 61: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_sample_completed_
      -- 
    ack_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1997_final_reg_ack_0, ack => convTransposeB_CP_4543_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_update_completed_
      -- 
    ack_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1997_final_reg_ack_1, ack => convTransposeB_CP_4543_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/ptr_deref_2000_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/ptr_deref_2000_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/ptr_deref_2000_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/ptr_deref_2000_Split/$entry
      -- 
    rr_5105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(63), ack => ptr_deref_2000_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(57) & convTransposeB_CP_4543_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Sample/word_access_start/word_0/ra
      -- 
    ra_5106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_store_0_ack_0, ack => convTransposeB_CP_4543_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/word_access_complete/word_0/ca
      -- 
    ca_5117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_store_0_ack_1, ack => convTransposeB_CP_4543_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_sample_completed_
      -- 
    ra_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2005_inst_ack_0, ack => convTransposeB_CP_4543_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_update_completed_
      -- 
    ca_5131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2005_inst_ack_1, ack => convTransposeB_CP_4543_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1753/R_cmp_2019_place
      -- CP-element group 68: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017__exit__
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018__entry__
      -- CP-element group 68: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/$exit
      -- CP-element group 68: 	 branch_block_stmt_1753/if_stmt_2018_else_link/$entry
      -- 
    branch_req_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(68), ack => if_stmt_2018_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(52) & convTransposeB_CP_4543_elements(59) & convTransposeB_CP_4543_elements(65) & convTransposeB_CP_4543_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1753/merge_stmt_2024_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1753/if_stmt_2018_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1753/if_stmt_2018_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1753/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1753/merge_stmt_2024__exit__
      -- CP-element group 69: 	 branch_block_stmt_1753/assign_stmt_2030__entry__
      -- CP-element group 69: 	 branch_block_stmt_1753/assign_stmt_2030__exit__
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1753/assign_stmt_2030/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/assign_stmt_2030/$exit
      -- CP-element group 69: 	 branch_block_stmt_1753/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1753/merge_stmt_2024_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/merge_stmt_2024_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1753/merge_stmt_2024_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2018_branch_ack_1, ack => convTransposeB_CP_4543_elements(69)); -- 
    rr_5476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(69), ack => type_cast_2092_inst_req_0); -- 
    cr_5481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(69), ack => type_cast_2092_inst_req_1); -- 
    rr_5499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(69), ack => type_cast_2088_inst_req_0); -- 
    cr_5504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(69), ack => type_cast_2088_inst_req_1); -- 
    rr_5522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(69), ack => type_cast_2079_inst_req_0); -- 
    cr_5527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(69), ack => type_cast_2079_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1753/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1753/merge_stmt_2032_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1753/merge_stmt_2032__exit__
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068__entry__
      -- CP-element group 70: 	 branch_block_stmt_1753/if_stmt_2018_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1753/if_stmt_2018_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/$entry
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1753/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1753/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1753/merge_stmt_2032_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1753/merge_stmt_2032_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1753/merge_stmt_2032_PhiAck/dummy
      -- 
    else_choice_transition_5148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2018_branch_ack_0, ack => convTransposeB_CP_4543_elements(70)); -- 
    rr_5164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(70), ack => type_cast_2046_inst_req_0); -- 
    cr_5169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(70), ack => type_cast_2046_inst_req_1); -- 
    cr_5183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(70), ack => type_cast_2062_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Sample/ra
      -- 
    ra_5165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2046_inst_ack_0, ack => convTransposeB_CP_4543_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2046_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Sample/rr
      -- 
    ca_5170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2046_inst_ack_1, ack => convTransposeB_CP_4543_elements(72)); -- 
    rr_5178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(72), ack => type_cast_2062_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Sample/ra
      -- 
    ra_5179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2062_inst_ack_0, ack => convTransposeB_CP_4543_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1753/R_cmp117_2070_place
      -- CP-element group 74: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068__exit__
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069__entry__
      -- CP-element group 74: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/$exit
      -- CP-element group 74: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1753/assign_stmt_2038_to_assign_stmt_2068/type_cast_2062_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1753/if_stmt_2069_else_link/$entry
      -- 
    ca_5184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2062_inst_ack_1, ack => convTransposeB_CP_4543_elements(74)); -- 
    branch_req_5192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(74), ack => if_stmt_2069_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1753/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1753/merge_stmt_2103__exit__
      -- CP-element group 75: 	 branch_block_stmt_1753/assign_stmt_2108__entry__
      -- CP-element group 75: 	 branch_block_stmt_1753/if_stmt_2069_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1753/if_stmt_2069_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1753/assign_stmt_2108/$entry
      -- CP-element group 75: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1753/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1753/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1753/merge_stmt_2103_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1753/merge_stmt_2103_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1753/merge_stmt_2103_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1753/merge_stmt_2103_PhiAck/dummy
      -- 
    if_choice_transition_5197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2069_branch_ack_1, ack => convTransposeB_CP_4543_elements(75)); -- 
    req_5217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(75), ack => WPIPE_Block1_done_2105_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	111 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/if_stmt_2069_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1753/if_stmt_2069_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2076/$entry
      -- CP-element group 76: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/$entry
      -- 
    else_choice_transition_5201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2069_branch_ack_0, ack => convTransposeB_CP_4543_elements(76)); -- 
    rr_5419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(76), ack => type_cast_2094_inst_req_0); -- 
    cr_5424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(76), ack => type_cast_2094_inst_req_1); -- 
    rr_5442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(76), ack => type_cast_2086_inst_req_0); -- 
    cr_5447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(76), ack => type_cast_2086_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Update/req
      -- 
    ack_5218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2105_inst_ack_0, ack => convTransposeB_CP_4543_elements(77)); -- 
    req_5222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(77), ack => WPIPE_Block1_done_2105_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1753/$exit
      -- CP-element group 78: 	 branch_block_stmt_1753/branch_block_stmt_1753__exit__
      -- CP-element group 78: 	 branch_block_stmt_1753/assign_stmt_2108__exit__
      -- CP-element group 78: 	 branch_block_stmt_1753/return__
      -- CP-element group 78: 	 branch_block_stmt_1753/merge_stmt_2110__exit__
      -- CP-element group 78: 	 branch_block_stmt_1753/assign_stmt_2108/$exit
      -- CP-element group 78: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1753/assign_stmt_2108/WPIPE_Block1_done_2105_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1753/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1753/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1753/merge_stmt_2110_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1753/merge_stmt_2110_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1753/merge_stmt_2110_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1753/merge_stmt_2110_PhiAck/dummy
      -- 
    ack_5223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2105_inst_ack_1, ack => convTransposeB_CP_4543_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Sample/ra
      -- 
    ra_5243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1892_inst_ack_0, ack => convTransposeB_CP_4543_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/Update/ca
      -- 
    ca_5248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1892_inst_ack_1, ack => convTransposeB_CP_4543_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/$exit
      -- CP-element group 81: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/$exit
      -- CP-element group 81: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1892/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_req
      -- 
    phi_stmt_1889_req_5249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1889_req_5249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(81), ack => phi_stmt_1889_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(79) & convTransposeB_CP_4543_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1882/$exit
      -- CP-element group 82: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1886_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_req
      -- 
    phi_stmt_1882_req_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1882_req_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(82), ack => phi_stmt_1882_req_0); -- 
    -- Element group convTransposeB_CP_4543_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4543_elements(43), ack => convTransposeB_CP_4543_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1875/$exit
      -- CP-element group 83: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1879_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_req
      -- 
    phi_stmt_1875_req_5265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1875_req_5265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(83), ack => phi_stmt_1875_req_0); -- 
    -- Element group convTransposeB_CP_4543_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4543_elements(43), ack => convTransposeB_CP_4543_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1868/$exit
      -- CP-element group 84: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1872_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_req
      -- 
    phi_stmt_1868_req_5273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_req_5273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(84), ack => phi_stmt_1868_req_0); -- 
    -- Element group convTransposeB_CP_4543_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4543_elements(43), ack => convTransposeB_CP_4543_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1753/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(81) & convTransposeB_CP_4543_elements(82) & convTransposeB_CP_4543_elements(83) & convTransposeB_CP_4543_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Sample/ra
      -- 
    ra_5293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_0, ack => convTransposeB_CP_4543_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/Update/ca
      -- 
    ca_5298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_1, ack => convTransposeB_CP_4543_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/$exit
      -- CP-element group 88: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/$exit
      -- CP-element group 88: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_sources/type_cast_1894/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1889/phi_stmt_1889_req
      -- 
    phi_stmt_1889_req_5299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1889_req_5299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(88), ack => phi_stmt_1889_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(86) & convTransposeB_CP_4543_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Sample/ra
      -- 
    ra_5316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_0, ack => convTransposeB_CP_4543_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/Update/ca
      -- 
    ca_5321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_1, ack => convTransposeB_CP_4543_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/$exit
      -- CP-element group 91: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/$exit
      -- CP-element group 91: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_sources/type_cast_1888/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1882/phi_stmt_1882_req
      -- 
    phi_stmt_1882_req_5322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1882_req_5322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(91), ack => phi_stmt_1882_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(89) & convTransposeB_CP_4543_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Sample/ra
      -- 
    ra_5339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_0, ack => convTransposeB_CP_4543_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/Update/ca
      -- 
    ca_5344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_1, ack => convTransposeB_CP_4543_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/$exit
      -- CP-element group 94: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/$exit
      -- CP-element group 94: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_sources/type_cast_1881/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1875/phi_stmt_1875_req
      -- 
    phi_stmt_1875_req_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1875_req_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(94), ack => phi_stmt_1875_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(92) & convTransposeB_CP_4543_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Sample/ra
      -- 
    ra_5362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1874_inst_ack_0, ack => convTransposeB_CP_4543_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/Update/ca
      -- 
    ca_5367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1874_inst_ack_1, ack => convTransposeB_CP_4543_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/$exit
      -- CP-element group 97: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/$exit
      -- CP-element group 97: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1868/phi_stmt_1868_req
      -- 
    phi_stmt_1868_req_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_req_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(97), ack => phi_stmt_1868_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(95) & convTransposeB_CP_4543_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1753/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(88) & convTransposeB_CP_4543_elements(91) & convTransposeB_CP_4543_elements(94) & convTransposeB_CP_4543_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1753/merge_stmt_1867_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1753/merge_stmt_1867_PhiAck/$entry
      -- 
    convTransposeB_CP_4543_elements(99) <= OrReduce(convTransposeB_CP_4543_elements(85) & convTransposeB_CP_4543_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1753/merge_stmt_1867_PhiAck/phi_stmt_1868_ack
      -- 
    phi_stmt_1868_ack_5373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1868_ack_0, ack => convTransposeB_CP_4543_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1753/merge_stmt_1867_PhiAck/phi_stmt_1875_ack
      -- 
    phi_stmt_1875_ack_5374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1875_ack_0, ack => convTransposeB_CP_4543_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1753/merge_stmt_1867_PhiAck/phi_stmt_1882_ack
      -- 
    phi_stmt_1882_ack_5375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1882_ack_0, ack => convTransposeB_CP_4543_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1753/merge_stmt_1867_PhiAck/phi_stmt_1889_ack
      -- 
    phi_stmt_1889_ack_5376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1889_ack_0, ack => convTransposeB_CP_4543_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_2000_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1996_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1753/merge_stmt_1867__exit__
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017__entry__
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1929_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1933_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1937_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_1967_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/type_cast_2005_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/array_obj_ref_1973_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1974_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/ptr_deref_1978_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1753/assign_stmt_1901_to_assign_stmt_2017/addr_of_1997_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1753/merge_stmt_1867_PhiAck/$exit
      -- 
    rr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_2005_inst_req_0); -- 
    cr_5116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => ptr_deref_2000_store_0_req_1); -- 
    req_5051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => array_obj_ref_1996_index_offset_req_1); -- 
    req_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => addr_of_1997_final_reg_req_1); -- 
    rr_4877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1929_inst_req_0); -- 
    cr_4882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1929_inst_req_1); -- 
    rr_4891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1933_inst_req_0); -- 
    cr_4896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1933_inst_req_1); -- 
    rr_4905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1937_inst_req_0); -- 
    cr_4910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1937_inst_req_1); -- 
    rr_4919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1967_inst_req_0); -- 
    cr_4924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_1967_inst_req_1); -- 
    cr_5130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => type_cast_2005_inst_req_1); -- 
    req_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => array_obj_ref_1973_index_offset_req_1); -- 
    req_4970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => addr_of_1974_final_reg_req_1); -- 
    cr_5015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(104), ack => ptr_deref_1978_load_0_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(100) & convTransposeB_CP_4543_elements(101) & convTransposeB_CP_4543_elements(102) & convTransposeB_CP_4543_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Sample/ra
      -- 
    ra_5420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2094_inst_ack_0, ack => convTransposeB_CP_4543_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/Update/ca
      -- 
    ca_5425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2094_inst_ack_1, ack => convTransposeB_CP_4543_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/$exit
      -- CP-element group 107: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/$exit
      -- CP-element group 107: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2094/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_req
      -- 
    phi_stmt_2089_req_5426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2089_req_5426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(107), ack => phi_stmt_2089_req_1); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(105) & convTransposeB_CP_4543_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/ra
      -- 
    ra_5443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2086_inst_ack_0, ack => convTransposeB_CP_4543_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/ca
      -- 
    ca_5448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2086_inst_ack_1, ack => convTransposeB_CP_4543_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/$exit
      -- CP-element group 110: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$exit
      -- CP-element group 110: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/$exit
      -- CP-element group 110: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/$exit
      -- CP-element group 110: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_req
      -- 
    phi_stmt_2083_req_5449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2083_req_5449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(110), ack => phi_stmt_2083_req_0); -- 
    convTransposeB_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(108) & convTransposeB_CP_4543_elements(109);
      gj_convTransposeB_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  output  delay-element  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	76 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2076/$exit
      -- CP-element group 111: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2082_konst_delay_trans
      -- CP-element group 111: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_req
      -- 
    phi_stmt_2076_req_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2076_req_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(111), ack => phi_stmt_2076_req_1); -- 
    -- Element group convTransposeB_CP_4543_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => convTransposeB_CP_4543_elements(76), ack => convTransposeB_CP_4543_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1753/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(107) & convTransposeB_CP_4543_elements(110) & convTransposeB_CP_4543_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Sample/ra
      -- 
    ra_5477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2092_inst_ack_0, ack => convTransposeB_CP_4543_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/Update/ca
      -- 
    ca_5482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2092_inst_ack_1, ack => convTransposeB_CP_4543_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/$exit
      -- CP-element group 115: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/$exit
      -- CP-element group 115: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_sources/type_cast_2092/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2089/phi_stmt_2089_req
      -- 
    phi_stmt_2089_req_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2089_req_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(115), ack => phi_stmt_2089_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(113) & convTransposeB_CP_4543_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Sample/ra
      -- 
    ra_5500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2088_inst_ack_0, ack => convTransposeB_CP_4543_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/Update/ca
      -- 
    ca_5505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2088_inst_ack_1, ack => convTransposeB_CP_4543_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/$exit
      -- CP-element group 118: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/$exit
      -- CP-element group 118: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2088/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2083/phi_stmt_2083_req
      -- 
    phi_stmt_2083_req_5506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2083_req_5506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(118), ack => phi_stmt_2083_req_1); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(116) & convTransposeB_CP_4543_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Sample/ra
      -- 
    ra_5523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2079_inst_ack_0, ack => convTransposeB_CP_4543_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/Update/ca
      -- 
    ca_5528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2079_inst_ack_1, ack => convTransposeB_CP_4543_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/$exit
      -- CP-element group 121: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/$exit
      -- CP-element group 121: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_sources/type_cast_2079/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2076/phi_stmt_2076_req
      -- 
    phi_stmt_2076_req_5529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2076_req_5529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4543_elements(121), ack => phi_stmt_2076_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(119) & convTransposeB_CP_4543_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1753/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(115) & convTransposeB_CP_4543_elements(118) & convTransposeB_CP_4543_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1753/merge_stmt_2075_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1753/merge_stmt_2075_PhiAck/$entry
      -- 
    convTransposeB_CP_4543_elements(123) <= OrReduce(convTransposeB_CP_4543_elements(112) & convTransposeB_CP_4543_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1753/merge_stmt_2075_PhiAck/phi_stmt_2076_ack
      -- 
    phi_stmt_2076_ack_5534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2076_ack_0, ack => convTransposeB_CP_4543_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1753/merge_stmt_2075_PhiAck/phi_stmt_2083_ack
      -- 
    phi_stmt_2083_ack_5535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2083_ack_0, ack => convTransposeB_CP_4543_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1753/merge_stmt_2075_PhiAck/phi_stmt_2089_ack
      -- 
    phi_stmt_2089_ack_5536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2089_ack_0, ack => convTransposeB_CP_4543_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1753/merge_stmt_2075_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4543_elements(124) & convTransposeB_CP_4543_elements(125) & convTransposeB_CP_4543_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4543_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_1995_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_1995_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1972_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1972_scaled : std_logic_vector(13 downto 0);
    signal add45_1827 : std_logic_vector(15 downto 0);
    signal add58_1838 : std_logic_vector(15 downto 0);
    signal add77_1948 : std_logic_vector(63 downto 0);
    signal add79_1958 : std_logic_vector(63 downto 0);
    signal add91_2012 : std_logic_vector(31 downto 0);
    signal add98_2030 : std_logic_vector(15 downto 0);
    signal add_1805 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1906 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1973_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1973_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1973_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1973_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1973_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1973_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1996_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1996_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1996_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1996_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1996_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1996_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_1975 : std_logic_vector(31 downto 0);
    signal arrayidx87_1998 : std_logic_vector(31 downto 0);
    signal call11_1774 : std_logic_vector(15 downto 0);
    signal call13_1777 : std_logic_vector(15 downto 0);
    signal call14_1780 : std_logic_vector(15 downto 0);
    signal call15_1783 : std_logic_vector(15 downto 0);
    signal call16_1796 : std_logic_vector(15 downto 0);
    signal call18_1808 : std_logic_vector(15 downto 0);
    signal call1_1759 : std_logic_vector(15 downto 0);
    signal call20_1811 : std_logic_vector(15 downto 0);
    signal call22_1814 : std_logic_vector(15 downto 0);
    signal call3_1762 : std_logic_vector(15 downto 0);
    signal call5_1765 : std_logic_vector(15 downto 0);
    signal call7_1768 : std_logic_vector(15 downto 0);
    signal call9_1771 : std_logic_vector(15 downto 0);
    signal call_1756 : std_logic_vector(15 downto 0);
    signal cmp106_2043 : std_logic_vector(0 downto 0);
    signal cmp117_2068 : std_logic_vector(0 downto 0);
    signal cmp_2017 : std_logic_vector(0 downto 0);
    signal conv112_2063 : std_logic_vector(31 downto 0);
    signal conv115_1859 : std_logic_vector(31 downto 0);
    signal conv17_1800 : std_logic_vector(31 downto 0);
    signal conv65_1930 : std_logic_vector(63 downto 0);
    signal conv68_1847 : std_logic_vector(63 downto 0);
    signal conv70_1934 : std_logic_vector(63 downto 0);
    signal conv73_1851 : std_logic_vector(63 downto 0);
    signal conv75_1938 : std_logic_vector(63 downto 0);
    signal conv90_2006 : std_logic_vector(31 downto 0);
    signal conv94_1855 : std_logic_vector(31 downto 0);
    signal conv_1787 : std_logic_vector(31 downto 0);
    signal idxprom86_1991 : std_logic_vector(63 downto 0);
    signal idxprom_1968 : std_logic_vector(63 downto 0);
    signal inc110_2047 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2052 : std_logic_vector(15 downto 0);
    signal inc_2038 : std_logic_vector(15 downto 0);
    signal indvar_1868 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2101 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2089 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1889 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2083 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1882 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2059 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2076 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1875 : std_logic_vector(15 downto 0);
    signal mul54_1921 : std_logic_vector(15 downto 0);
    signal mul76_1943 : std_logic_vector(63 downto 0);
    signal mul78_1953 : std_logic_vector(63 downto 0);
    signal mul_1911 : std_logic_vector(15 downto 0);
    signal ptr_deref_1978_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1978_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1978_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1978_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1978_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2000_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2000_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2000_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2000_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2000_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2000_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1793 : std_logic_vector(31 downto 0);
    signal shr116132_1865 : std_logic_vector(31 downto 0);
    signal shr131_1821 : std_logic_vector(15 downto 0);
    signal shr81_1964 : std_logic_vector(31 downto 0);
    signal shr85_1985 : std_logic_vector(63 downto 0);
    signal sub48_1916 : std_logic_vector(15 downto 0);
    signal sub61_1843 : std_logic_vector(15 downto 0);
    signal sub62_1926 : std_logic_vector(15 downto 0);
    signal sub_1832 : std_logic_vector(15 downto 0);
    signal tmp1_1901 : std_logic_vector(31 downto 0);
    signal tmp83_1979 : std_logic_vector(63 downto 0);
    signal type_cast_1791_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1819_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1825_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1836_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1863_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1872_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1874_wire : std_logic_vector(31 downto 0);
    signal type_cast_1879_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1881_wire : std_logic_vector(15 downto 0);
    signal type_cast_1886_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1888_wire : std_logic_vector(15 downto 0);
    signal type_cast_1892_wire : std_logic_vector(15 downto 0);
    signal type_cast_1894_wire : std_logic_vector(15 downto 0);
    signal type_cast_1899_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1983_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1989_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2010_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2028_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2036_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2056_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2079_wire : std_logic_vector(15 downto 0);
    signal type_cast_2082_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2086_wire : std_logic_vector(15 downto 0);
    signal type_cast_2088_wire : std_logic_vector(15 downto 0);
    signal type_cast_2092_wire : std_logic_vector(15 downto 0);
    signal type_cast_2094_wire : std_logic_vector(15 downto 0);
    signal type_cast_2099_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2107_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1973_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1973_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1973_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1973_resized_base_address <= "00000000000000";
    array_obj_ref_1996_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1996_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1996_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1996_resized_base_address <= "00000000000000";
    ptr_deref_1978_word_offset_0 <= "00000000000000";
    ptr_deref_2000_word_offset_0 <= "00000000000000";
    type_cast_1791_wire_constant <= "00000000000000000000000000010000";
    type_cast_1819_wire_constant <= "0000000000000010";
    type_cast_1825_wire_constant <= "1111111111111111";
    type_cast_1836_wire_constant <= "1111111111111111";
    type_cast_1863_wire_constant <= "00000000000000000000000000000001";
    type_cast_1872_wire_constant <= "00000000000000000000000000000000";
    type_cast_1879_wire_constant <= "0000000000000000";
    type_cast_1886_wire_constant <= "0000000000000000";
    type_cast_1899_wire_constant <= "00000000000000000000000000000100";
    type_cast_1962_wire_constant <= "00000000000000000000000000000010";
    type_cast_1983_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1989_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2010_wire_constant <= "00000000000000000000000000000100";
    type_cast_2028_wire_constant <= "0000000000000100";
    type_cast_2036_wire_constant <= "0000000000000001";
    type_cast_2056_wire_constant <= "0000000000000000";
    type_cast_2082_wire_constant <= "0000000000000000";
    type_cast_2099_wire_constant <= "00000000000000000000000000000001";
    type_cast_2107_wire_constant <= "0000000000000001";
    phi_stmt_1868: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1872_wire_constant & type_cast_1874_wire;
      req <= phi_stmt_1868_req_0 & phi_stmt_1868_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1868",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1868_ack_0,
          idata => idata,
          odata => indvar_1868,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1868
    phi_stmt_1875: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1879_wire_constant & type_cast_1881_wire;
      req <= phi_stmt_1875_req_0 & phi_stmt_1875_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1875",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1875_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1875,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1875
    phi_stmt_1882: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1886_wire_constant & type_cast_1888_wire;
      req <= phi_stmt_1882_req_0 & phi_stmt_1882_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1882",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1882_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1882,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1882
    phi_stmt_1889: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1892_wire & type_cast_1894_wire;
      req <= phi_stmt_1889_req_0 & phi_stmt_1889_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1889",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1889_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1889,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1889
    phi_stmt_2076: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2079_wire & type_cast_2082_wire_constant;
      req <= phi_stmt_2076_req_0 & phi_stmt_2076_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2076",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2076_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2076,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2076
    phi_stmt_2083: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2086_wire & type_cast_2088_wire;
      req <= phi_stmt_2083_req_0 & phi_stmt_2083_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2083",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2083_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2083,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2083
    phi_stmt_2089: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2092_wire & type_cast_2094_wire;
      req <= phi_stmt_2089_req_0 & phi_stmt_2089_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2089",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2089_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2089,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2089
    -- flow-through select operator MUX_2058_inst
    input_dim1x_x2_2059 <= type_cast_2056_wire_constant when (cmp106_2043(0) /=  '0') else inc_2038;
    addr_of_1974_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1974_final_reg_req_0;
      addr_of_1974_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1974_final_reg_req_1;
      addr_of_1974_final_reg_ack_1<= rack(0);
      addr_of_1974_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1974_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1973_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1975,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1997_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1997_final_reg_req_0;
      addr_of_1997_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1997_final_reg_req_1;
      addr_of_1997_final_reg_ack_1<= rack(0);
      addr_of_1997_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1997_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1996_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_1998,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1786_inst_req_0;
      type_cast_1786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1786_inst_req_1;
      type_cast_1786_inst_ack_1<= rack(0);
      type_cast_1786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1799_inst_req_0;
      type_cast_1799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1799_inst_req_1;
      type_cast_1799_inst_ack_1<= rack(0);
      type_cast_1799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1846_inst_req_0;
      type_cast_1846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1846_inst_req_1;
      type_cast_1846_inst_ack_1<= rack(0);
      type_cast_1846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1847,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1850_inst_req_0;
      type_cast_1850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1850_inst_req_1;
      type_cast_1850_inst_ack_1<= rack(0);
      type_cast_1850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1854_inst_req_0;
      type_cast_1854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1854_inst_req_1;
      type_cast_1854_inst_ack_1<= rack(0);
      type_cast_1854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1762,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1858_inst_req_0;
      type_cast_1858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1858_inst_req_1;
      type_cast_1858_inst_ack_1<= rack(0);
      type_cast_1858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1874_inst_req_0;
      type_cast_1874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1874_inst_req_1;
      type_cast_1874_inst_ack_1<= rack(0);
      type_cast_1874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1874_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1881_inst_req_0;
      type_cast_1881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1881_inst_req_1;
      type_cast_1881_inst_ack_1<= rack(0);
      type_cast_1881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2076,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1881_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1888_inst_req_0;
      type_cast_1888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1888_inst_req_1;
      type_cast_1888_inst_ack_1<= rack(0);
      type_cast_1888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1888_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1888_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1892_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1892_inst_req_0;
      type_cast_1892_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1892_inst_req_1;
      type_cast_1892_inst_ack_1<= rack(0);
      type_cast_1892_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1892_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1892_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1894_inst_req_0;
      type_cast_1894_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1894_inst_req_1;
      type_cast_1894_inst_ack_1<= rack(0);
      type_cast_1894_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1894_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2089,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1894_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1929_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1929_inst_req_0;
      type_cast_1929_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1929_inst_req_1;
      type_cast_1929_inst_ack_1<= rack(0);
      type_cast_1929_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1929_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_1930,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1933_inst_req_0;
      type_cast_1933_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1933_inst_req_1;
      type_cast_1933_inst_ack_1<= rack(0);
      type_cast_1933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_1926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1937_inst_req_0;
      type_cast_1937_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1937_inst_req_1;
      type_cast_1937_inst_ack_1<= rack(0);
      type_cast_1937_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1937_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_1916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1938,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1967_inst_req_0;
      type_cast_1967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1967_inst_req_1;
      type_cast_1967_inst_ack_1<= rack(0);
      type_cast_1967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_1964,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2005_inst_req_0;
      type_cast_2005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2005_inst_req_1;
      type_cast_2005_inst_ack_1<= rack(0);
      type_cast_2005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2006,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2046_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2046_inst_req_0;
      type_cast_2046_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2046_inst_req_1;
      type_cast_2046_inst_ack_1<= rack(0);
      type_cast_2046_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2046_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2043,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2047,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2062_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2062_inst_req_0;
      type_cast_2062_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2062_inst_req_1;
      type_cast_2062_inst_ack_1<= rack(0);
      type_cast_2062_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2062_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2063,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2079_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2079_inst_req_0;
      type_cast_2079_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2079_inst_req_1;
      type_cast_2079_inst_ack_1<= rack(0);
      type_cast_2079_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2079_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2079_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2086_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2086_inst_req_0;
      type_cast_2086_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2086_inst_req_1;
      type_cast_2086_inst_ack_1<= rack(0);
      type_cast_2086_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2086_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2059,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2086_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2088_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2088_inst_req_0;
      type_cast_2088_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2088_inst_req_1;
      type_cast_2088_inst_ack_1<= rack(0);
      type_cast_2088_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2088_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2088_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2092_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2092_inst_req_0;
      type_cast_2092_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2092_inst_req_1;
      type_cast_2092_inst_ack_1<= rack(0);
      type_cast_2092_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2092_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2092_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2094_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2094_inst_req_0;
      type_cast_2094_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2094_inst_req_1;
      type_cast_2094_inst_ack_1<= rack(0);
      type_cast_2094_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2094_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2094_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1973_index_1_rename
    process(R_idxprom_1972_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1972_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1972_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1973_index_1_resize
    process(idxprom_1968) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1968;
      ov := iv(13 downto 0);
      R_idxprom_1972_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1973_root_address_inst
    process(array_obj_ref_1973_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1973_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1973_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1996_index_1_rename
    process(R_idxprom86_1995_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_1995_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_1995_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1996_index_1_resize
    process(idxprom86_1991) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_1991;
      ov := iv(13 downto 0);
      R_idxprom86_1995_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1996_root_address_inst
    process(array_obj_ref_1996_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1996_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1996_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1978_addr_0
    process(ptr_deref_1978_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1978_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1978_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1978_base_resize
    process(arrayidx82_1975) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1975;
      ov := iv(13 downto 0);
      ptr_deref_1978_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1978_gather_scatter
    process(ptr_deref_1978_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1978_data_0;
      ov(63 downto 0) := iv;
      tmp83_1979 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1978_root_address_inst
    process(ptr_deref_1978_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1978_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1978_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2000_addr_0
    process(ptr_deref_2000_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2000_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2000_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2000_base_resize
    process(arrayidx87_1998) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_1998;
      ov := iv(13 downto 0);
      ptr_deref_2000_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2000_gather_scatter
    process(tmp83_1979) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_1979;
      ov(63 downto 0) := iv;
      ptr_deref_2000_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2000_root_address_inst
    process(ptr_deref_2000_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2000_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2000_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2018_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2017;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2018_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2018_branch_req_0,
          ack0 => if_stmt_2018_branch_ack_0,
          ack1 => if_stmt_2018_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2069_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2068;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2069_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2069_branch_req_0,
          ack0 => if_stmt_2069_branch_ack_0,
          ack1 => if_stmt_2069_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1826_inst
    process(call7_1768) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1768, type_cast_1825_wire_constant, tmp_var);
      add45_1827 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1837_inst
    process(call9_1771) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1771, type_cast_1836_wire_constant, tmp_var);
      add58_1838 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1915_inst
    process(sub_1832, mul_1911) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1832, mul_1911, tmp_var);
      sub48_1916 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1925_inst
    process(sub61_1843, mul54_1921) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1843, mul54_1921, tmp_var);
      sub62_1926 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2029_inst
    process(input_dim2x_x1_1875) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1875, type_cast_2028_wire_constant, tmp_var);
      add98_2030 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2037_inst
    process(input_dim1x_x1_1882) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1882, type_cast_2036_wire_constant, tmp_var);
      inc_2038 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2051_inst
    process(inc110_2047, input_dim0x_x2_1889) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2047, input_dim0x_x2_1889, tmp_var);
      inc110x_xinput_dim0x_x2_2052 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1905_inst
    process(add_1805, tmp1_1901) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1805, tmp1_1901, tmp_var);
      add_src_0x_x0_1906 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2011_inst
    process(conv90_2006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2006, type_cast_2010_wire_constant, tmp_var);
      add91_2012 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2100_inst
    process(indvar_1868) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1868, type_cast_2099_wire_constant, tmp_var);
      indvarx_xnext_2101 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1947_inst
    process(mul76_1943, conv70_1934) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_1943, conv70_1934, tmp_var);
      add77_1948 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1957_inst
    process(mul78_1953, conv65_1930) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_1953, conv65_1930, tmp_var);
      add79_1958 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1990_inst
    process(shr85_1985) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_1985, type_cast_1989_wire_constant, tmp_var);
      idxprom86_1991 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2042_inst
    process(inc_2038, call1_1759) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2038, call1_1759, tmp_var);
      cmp106_2043 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2067_inst
    process(conv112_2063, shr116132_1865) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2063, shr116132_1865, tmp_var);
      cmp117_2068 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1820_inst
    process(call_1756) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1756, type_cast_1819_wire_constant, tmp_var);
      shr131_1821 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1864_inst
    process(conv115_1859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1859, type_cast_1863_wire_constant, tmp_var);
      shr116132_1865 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1963_inst
    process(add_src_0x_x0_1906) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1906, type_cast_1962_wire_constant, tmp_var);
      shr81_1964 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1984_inst
    process(add79_1958) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_1958, type_cast_1983_wire_constant, tmp_var);
      shr85_1985 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1910_inst
    process(input_dim0x_x2_1889, call13_1777) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1889, call13_1777, tmp_var);
      mul_1911 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1920_inst
    process(input_dim1x_x1_1882, call13_1777) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1882, call13_1777, tmp_var);
      mul54_1921 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1900_inst
    process(indvar_1868) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1868, type_cast_1899_wire_constant, tmp_var);
      tmp1_1901 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1942_inst
    process(conv75_1938, conv73_1851) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_1938, conv73_1851, tmp_var);
      mul76_1943 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1952_inst
    process(add77_1948, conv68_1847) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_1948, conv68_1847, tmp_var);
      mul78_1953 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1804_inst
    process(shl_1793, conv17_1800) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1793, conv17_1800, tmp_var);
      add_1805 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1792_inst
    process(conv_1787) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1787, type_cast_1791_wire_constant, tmp_var);
      shl_1793 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1831_inst
    process(add45_1827, call14_1780) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1827, call14_1780, tmp_var);
      sub_1832 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1842_inst
    process(add58_1838, call14_1780) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1838, call14_1780, tmp_var);
      sub61_1843 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2016_inst
    process(add91_2012, conv94_1855) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2012, conv94_1855, tmp_var);
      cmp_2017 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_1973_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1972_scaled;
      array_obj_ref_1973_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1973_index_offset_req_0;
      array_obj_ref_1973_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1973_index_offset_req_1;
      array_obj_ref_1973_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_1996_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_1995_scaled;
      array_obj_ref_1996_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1996_index_offset_req_0;
      array_obj_ref_1996_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1996_index_offset_req_1;
      array_obj_ref_1996_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_1978_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1978_load_0_req_0;
      ptr_deref_1978_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1978_load_0_req_1;
      ptr_deref_1978_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1978_word_address_0;
      ptr_deref_1978_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2000_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2000_store_0_req_0;
      ptr_deref_2000_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2000_store_0_req_1;
      ptr_deref_2000_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2000_word_address_0;
      data_in <= ptr_deref_2000_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1755_inst RPIPE_Block1_start_1758_inst RPIPE_Block1_start_1761_inst RPIPE_Block1_start_1764_inst RPIPE_Block1_start_1767_inst RPIPE_Block1_start_1770_inst RPIPE_Block1_start_1773_inst RPIPE_Block1_start_1776_inst RPIPE_Block1_start_1779_inst RPIPE_Block1_start_1782_inst RPIPE_Block1_start_1795_inst RPIPE_Block1_start_1807_inst RPIPE_Block1_start_1810_inst RPIPE_Block1_start_1813_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1755_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1758_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1761_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1764_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1767_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1770_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1773_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1776_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1779_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1782_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1795_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1807_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1810_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1813_inst_req_0;
      RPIPE_Block1_start_1755_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1758_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1761_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1764_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1767_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1770_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1773_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1776_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1779_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1782_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1795_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1807_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1810_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1813_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1755_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1758_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1761_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1764_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1767_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1770_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1773_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1776_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1779_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1782_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1795_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1807_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1810_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1813_inst_req_1;
      RPIPE_Block1_start_1755_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1758_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1761_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1764_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1767_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1770_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1773_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1776_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1779_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1782_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1795_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1807_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1810_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1813_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_1756 <= data_out(223 downto 208);
      call1_1759 <= data_out(207 downto 192);
      call3_1762 <= data_out(191 downto 176);
      call5_1765 <= data_out(175 downto 160);
      call7_1768 <= data_out(159 downto 144);
      call9_1771 <= data_out(143 downto 128);
      call11_1774 <= data_out(127 downto 112);
      call13_1777 <= data_out(111 downto 96);
      call14_1780 <= data_out(95 downto 80);
      call15_1783 <= data_out(79 downto 64);
      call16_1796 <= data_out(63 downto 48);
      call18_1808 <= data_out(47 downto 32);
      call20_1811 <= data_out(31 downto 16);
      call22_1814 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2105_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2105_inst_req_0;
      WPIPE_Block1_done_2105_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2105_inst_req_1;
      WPIPE_Block1_done_2105_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2107_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5553_start: Boolean;
  signal convTransposeC_CP_5553_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2418_inst_req_1 : boolean;
  signal addr_of_2369_final_reg_ack_0 : boolean;
  signal RPIPE_Block2_start_2116_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2116_inst_ack_1 : boolean;
  signal if_stmt_2390_branch_ack_0 : boolean;
  signal addr_of_2369_final_reg_req_0 : boolean;
  signal RPIPE_Block2_start_2116_inst_ack_0 : boolean;
  signal type_cast_2418_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2116_inst_req_0 : boolean;
  signal addr_of_2369_final_reg_req_1 : boolean;
  signal if_stmt_2390_branch_ack_1 : boolean;
  signal RPIPE_Block2_start_2122_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2122_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2119_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2119_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2119_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2119_inst_req_0 : boolean;
  signal ptr_deref_2372_store_0_req_0 : boolean;
  signal addr_of_2369_final_reg_ack_1 : boolean;
  signal ptr_deref_2372_store_0_ack_0 : boolean;
  signal type_cast_2434_inst_req_1 : boolean;
  signal type_cast_2434_inst_ack_1 : boolean;
  signal if_stmt_2441_branch_ack_1 : boolean;
  signal type_cast_2434_inst_req_0 : boolean;
  signal if_stmt_2390_branch_req_0 : boolean;
  signal type_cast_2434_inst_ack_0 : boolean;
  signal ptr_deref_2372_store_0_req_1 : boolean;
  signal ptr_deref_2372_store_0_ack_1 : boolean;
  signal type_cast_2377_inst_req_0 : boolean;
  signal if_stmt_2441_branch_req_0 : boolean;
  signal if_stmt_2441_branch_ack_0 : boolean;
  signal type_cast_2377_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2122_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2122_inst_ack_1 : boolean;
  signal array_obj_ref_2368_index_offset_ack_1 : boolean;
  signal array_obj_ref_2368_index_offset_req_1 : boolean;
  signal array_obj_ref_2368_index_offset_ack_0 : boolean;
  signal array_obj_ref_2368_index_offset_req_0 : boolean;
  signal RPIPE_Block2_start_2125_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2125_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2125_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2125_inst_ack_1 : boolean;
  signal type_cast_2377_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2128_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2128_inst_ack_0 : boolean;
  signal type_cast_2377_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2128_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2128_inst_ack_1 : boolean;
  signal type_cast_2418_inst_ack_0 : boolean;
  signal type_cast_2418_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2131_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2131_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2131_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2131_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2134_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2134_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2134_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2134_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2137_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2137_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2137_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2137_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2140_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2140_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2140_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2140_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2143_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2143_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2143_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2143_inst_ack_1 : boolean;
  signal type_cast_2147_inst_req_0 : boolean;
  signal type_cast_2147_inst_ack_0 : boolean;
  signal type_cast_2147_inst_req_1 : boolean;
  signal type_cast_2147_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2156_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2156_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2156_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2156_inst_ack_1 : boolean;
  signal type_cast_2160_inst_req_0 : boolean;
  signal type_cast_2160_inst_ack_0 : boolean;
  signal type_cast_2160_inst_req_1 : boolean;
  signal type_cast_2160_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2168_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2168_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2168_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2168_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2171_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2171_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2171_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2171_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2174_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2174_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2174_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2174_inst_ack_1 : boolean;
  signal type_cast_2207_inst_req_0 : boolean;
  signal type_cast_2207_inst_ack_0 : boolean;
  signal type_cast_2207_inst_req_1 : boolean;
  signal type_cast_2207_inst_ack_1 : boolean;
  signal type_cast_2211_inst_req_0 : boolean;
  signal type_cast_2211_inst_ack_0 : boolean;
  signal type_cast_2211_inst_req_1 : boolean;
  signal type_cast_2211_inst_ack_1 : boolean;
  signal type_cast_2215_inst_req_0 : boolean;
  signal type_cast_2215_inst_ack_0 : boolean;
  signal type_cast_2215_inst_req_1 : boolean;
  signal type_cast_2215_inst_ack_1 : boolean;
  signal type_cast_2219_inst_req_0 : boolean;
  signal type_cast_2219_inst_ack_0 : boolean;
  signal type_cast_2219_inst_req_1 : boolean;
  signal type_cast_2219_inst_ack_1 : boolean;
  signal type_cast_2301_inst_req_0 : boolean;
  signal type_cast_2301_inst_ack_0 : boolean;
  signal type_cast_2301_inst_req_1 : boolean;
  signal type_cast_2301_inst_ack_1 : boolean;
  signal type_cast_2305_inst_req_0 : boolean;
  signal type_cast_2305_inst_ack_0 : boolean;
  signal type_cast_2305_inst_req_1 : boolean;
  signal type_cast_2305_inst_ack_1 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal type_cast_2309_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_1 : boolean;
  signal type_cast_2339_inst_req_0 : boolean;
  signal type_cast_2339_inst_ack_0 : boolean;
  signal type_cast_2339_inst_req_1 : boolean;
  signal type_cast_2339_inst_ack_1 : boolean;
  signal array_obj_ref_2345_index_offset_req_0 : boolean;
  signal array_obj_ref_2345_index_offset_ack_0 : boolean;
  signal array_obj_ref_2345_index_offset_req_1 : boolean;
  signal array_obj_ref_2345_index_offset_ack_1 : boolean;
  signal addr_of_2346_final_reg_req_0 : boolean;
  signal addr_of_2346_final_reg_ack_0 : boolean;
  signal addr_of_2346_final_reg_req_1 : boolean;
  signal addr_of_2346_final_reg_ack_1 : boolean;
  signal ptr_deref_2350_load_0_req_0 : boolean;
  signal ptr_deref_2350_load_0_ack_0 : boolean;
  signal ptr_deref_2350_load_0_req_1 : boolean;
  signal ptr_deref_2350_load_0_ack_1 : boolean;
  signal WPIPE_Block2_done_2477_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2477_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2477_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2477_inst_ack_1 : boolean;
  signal phi_stmt_2240_req_0 : boolean;
  signal phi_stmt_2247_req_0 : boolean;
  signal type_cast_2266_inst_req_0 : boolean;
  signal type_cast_2266_inst_ack_0 : boolean;
  signal type_cast_2266_inst_req_1 : boolean;
  signal type_cast_2266_inst_ack_1 : boolean;
  signal phi_stmt_2261_req_1 : boolean;
  signal phi_stmt_2254_req_0 : boolean;
  signal type_cast_2246_inst_req_0 : boolean;
  signal type_cast_2246_inst_ack_0 : boolean;
  signal type_cast_2246_inst_req_1 : boolean;
  signal type_cast_2246_inst_ack_1 : boolean;
  signal phi_stmt_2240_req_1 : boolean;
  signal type_cast_2253_inst_req_0 : boolean;
  signal type_cast_2253_inst_ack_0 : boolean;
  signal type_cast_2253_inst_req_1 : boolean;
  signal type_cast_2253_inst_ack_1 : boolean;
  signal phi_stmt_2247_req_1 : boolean;
  signal type_cast_2264_inst_req_0 : boolean;
  signal type_cast_2264_inst_ack_0 : boolean;
  signal type_cast_2264_inst_req_1 : boolean;
  signal type_cast_2264_inst_ack_1 : boolean;
  signal phi_stmt_2261_req_0 : boolean;
  signal type_cast_2260_inst_req_0 : boolean;
  signal type_cast_2260_inst_ack_0 : boolean;
  signal type_cast_2260_inst_req_1 : boolean;
  signal type_cast_2260_inst_ack_1 : boolean;
  signal phi_stmt_2254_req_1 : boolean;
  signal phi_stmt_2240_ack_0 : boolean;
  signal phi_stmt_2247_ack_0 : boolean;
  signal phi_stmt_2254_ack_0 : boolean;
  signal phi_stmt_2261_ack_0 : boolean;
  signal phi_stmt_2448_req_0 : boolean;
  signal type_cast_2458_inst_req_0 : boolean;
  signal type_cast_2458_inst_ack_0 : boolean;
  signal type_cast_2458_inst_req_1 : boolean;
  signal type_cast_2458_inst_ack_1 : boolean;
  signal phi_stmt_2455_req_0 : boolean;
  signal type_cast_2464_inst_req_0 : boolean;
  signal type_cast_2464_inst_ack_0 : boolean;
  signal type_cast_2464_inst_req_1 : boolean;
  signal type_cast_2464_inst_ack_1 : boolean;
  signal phi_stmt_2461_req_0 : boolean;
  signal type_cast_2454_inst_req_0 : boolean;
  signal type_cast_2454_inst_ack_0 : boolean;
  signal type_cast_2454_inst_req_1 : boolean;
  signal type_cast_2454_inst_ack_1 : boolean;
  signal phi_stmt_2448_req_1 : boolean;
  signal type_cast_2460_inst_req_0 : boolean;
  signal type_cast_2460_inst_ack_0 : boolean;
  signal type_cast_2460_inst_req_1 : boolean;
  signal type_cast_2460_inst_ack_1 : boolean;
  signal phi_stmt_2455_req_1 : boolean;
  signal type_cast_2466_inst_req_0 : boolean;
  signal type_cast_2466_inst_ack_0 : boolean;
  signal type_cast_2466_inst_req_1 : boolean;
  signal type_cast_2466_inst_ack_1 : boolean;
  signal phi_stmt_2461_req_1 : boolean;
  signal phi_stmt_2448_ack_0 : boolean;
  signal phi_stmt_2455_ack_0 : boolean;
  signal phi_stmt_2461_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5553_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5553_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5553_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5553_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5553: Block -- control-path 
    signal convTransposeC_CP_5553_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5553_elements(0) <= convTransposeC_CP_5553_start;
    convTransposeC_CP_5553_symbol <= convTransposeC_CP_5553_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/$entry
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2114/$entry
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2114/branch_block_stmt_2114__entry__
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Update/cr
      -- 
    rr_5601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(0), ack => RPIPE_Block2_start_2116_inst_req_0); -- 
    cr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(0), ack => type_cast_2147_inst_req_1); -- 
    cr_5774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(0), ack => type_cast_2160_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2114/assign_stmt_2473__exit__
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2114/merge_stmt_2447__exit__
      -- CP-element group 1: 	 branch_block_stmt_2114/assign_stmt_2473__entry__
      -- CP-element group 1: 	 branch_block_stmt_2114/assign_stmt_2473/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/assign_stmt_2473/$exit
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Update/cr
      -- 
    rr_6302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2246_inst_req_0); -- 
    cr_6307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2246_inst_req_1); -- 
    rr_6325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2253_inst_req_0); -- 
    cr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2253_inst_req_1); -- 
    rr_6348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2264_inst_req_0); -- 
    cr_6353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2264_inst_req_1); -- 
    rr_6371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2260_inst_req_0); -- 
    cr_6376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(1), ack => type_cast_2260_inst_req_1); -- 
    convTransposeC_CP_5553_elements(1) <= convTransposeC_CP_5553_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Sample/$exit
      -- 
    ra_5602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2116_inst_ack_0, ack => convTransposeC_CP_5553_elements(2)); -- 
    cr_5606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(2), ack => RPIPE_Block2_start_2116_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2116_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Sample/$entry
      -- 
    ca_5607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2116_inst_ack_1, ack => convTransposeC_CP_5553_elements(3)); -- 
    rr_5615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(3), ack => RPIPE_Block2_start_2119_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Sample/$exit
      -- 
    ra_5616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2119_inst_ack_0, ack => convTransposeC_CP_5553_elements(4)); -- 
    cr_5620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(4), ack => RPIPE_Block2_start_2119_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2119_Update/$exit
      -- 
    ca_5621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2119_inst_ack_1, ack => convTransposeC_CP_5553_elements(5)); -- 
    rr_5629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(5), ack => RPIPE_Block2_start_2122_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Update/cr
      -- 
    ra_5630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2122_inst_ack_0, ack => convTransposeC_CP_5553_elements(6)); -- 
    cr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(6), ack => RPIPE_Block2_start_2122_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2122_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Sample/rr
      -- 
    ca_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2122_inst_ack_1, ack => convTransposeC_CP_5553_elements(7)); -- 
    rr_5643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(7), ack => RPIPE_Block2_start_2125_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Update/cr
      -- 
    ra_5644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2125_inst_ack_0, ack => convTransposeC_CP_5553_elements(8)); -- 
    cr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(8), ack => RPIPE_Block2_start_2125_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2125_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Sample/rr
      -- 
    ca_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2125_inst_ack_1, ack => convTransposeC_CP_5553_elements(9)); -- 
    rr_5657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(9), ack => RPIPE_Block2_start_2128_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Update/cr
      -- 
    ra_5658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2128_inst_ack_0, ack => convTransposeC_CP_5553_elements(10)); -- 
    cr_5662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(10), ack => RPIPE_Block2_start_2128_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2128_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Sample/rr
      -- 
    ca_5663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2128_inst_ack_1, ack => convTransposeC_CP_5553_elements(11)); -- 
    rr_5671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(11), ack => RPIPE_Block2_start_2131_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Update/cr
      -- 
    ra_5672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2131_inst_ack_0, ack => convTransposeC_CP_5553_elements(12)); -- 
    cr_5676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(12), ack => RPIPE_Block2_start_2131_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2131_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Sample/rr
      -- 
    ca_5677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2131_inst_ack_1, ack => convTransposeC_CP_5553_elements(13)); -- 
    rr_5685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(13), ack => RPIPE_Block2_start_2134_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Update/cr
      -- 
    ra_5686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2134_inst_ack_0, ack => convTransposeC_CP_5553_elements(14)); -- 
    cr_5690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(14), ack => RPIPE_Block2_start_2134_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2134_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Sample/rr
      -- 
    ca_5691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2134_inst_ack_1, ack => convTransposeC_CP_5553_elements(15)); -- 
    rr_5699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(15), ack => RPIPE_Block2_start_2137_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Update/cr
      -- 
    ra_5700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2137_inst_ack_0, ack => convTransposeC_CP_5553_elements(16)); -- 
    cr_5704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(16), ack => RPIPE_Block2_start_2137_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2137_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Sample/rr
      -- 
    ca_5705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2137_inst_ack_1, ack => convTransposeC_CP_5553_elements(17)); -- 
    rr_5713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(17), ack => RPIPE_Block2_start_2140_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Update/cr
      -- 
    ra_5714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2140_inst_ack_0, ack => convTransposeC_CP_5553_elements(18)); -- 
    cr_5718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(18), ack => RPIPE_Block2_start_2140_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2140_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Sample/rr
      -- 
    ca_5719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2140_inst_ack_1, ack => convTransposeC_CP_5553_elements(19)); -- 
    rr_5727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(19), ack => RPIPE_Block2_start_2143_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Update/cr
      -- 
    ra_5728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2143_inst_ack_0, ack => convTransposeC_CP_5553_elements(20)); -- 
    cr_5732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(20), ack => RPIPE_Block2_start_2143_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2143_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Sample/rr
      -- 
    ca_5733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2143_inst_ack_1, ack => convTransposeC_CP_5553_elements(21)); -- 
    rr_5741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(21), ack => type_cast_2147_inst_req_0); -- 
    rr_5755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(21), ack => RPIPE_Block2_start_2156_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Sample/ra
      -- 
    ra_5742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_0, ack => convTransposeC_CP_5553_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2147_Update/ca
      -- 
    ca_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_1, ack => convTransposeC_CP_5553_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Update/cr
      -- 
    ra_5756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2156_inst_ack_0, ack => convTransposeC_CP_5553_elements(24)); -- 
    cr_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(24), ack => RPIPE_Block2_start_2156_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2156_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Sample/rr
      -- 
    ca_5761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2156_inst_ack_1, ack => convTransposeC_CP_5553_elements(25)); -- 
    rr_5769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(25), ack => type_cast_2160_inst_req_0); -- 
    rr_5783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(25), ack => RPIPE_Block2_start_2168_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Sample/ra
      -- 
    ra_5770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2160_inst_ack_0, ack => convTransposeC_CP_5553_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/type_cast_2160_Update/ca
      -- 
    ca_5775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2160_inst_ack_1, ack => convTransposeC_CP_5553_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Update/cr
      -- 
    ra_5784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2168_inst_ack_0, ack => convTransposeC_CP_5553_elements(28)); -- 
    cr_5788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(28), ack => RPIPE_Block2_start_2168_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2168_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Sample/rr
      -- 
    ca_5789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2168_inst_ack_1, ack => convTransposeC_CP_5553_elements(29)); -- 
    rr_5797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(29), ack => RPIPE_Block2_start_2171_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Update/cr
      -- 
    ra_5798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2171_inst_ack_0, ack => convTransposeC_CP_5553_elements(30)); -- 
    cr_5802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(30), ack => RPIPE_Block2_start_2171_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2171_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Sample/rr
      -- 
    ca_5803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2171_inst_ack_1, ack => convTransposeC_CP_5553_elements(31)); -- 
    rr_5811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(31), ack => RPIPE_Block2_start_2174_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Update/cr
      -- 
    ra_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2174_inst_ack_0, ack => convTransposeC_CP_5553_elements(32)); -- 
    cr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(32), ack => RPIPE_Block2_start_2174_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/RPIPE_Block2_start_2174_Update/ca
      -- 
    ca_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2174_inst_ack_1, ack => convTransposeC_CP_5553_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175/$exit
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2117_to_assign_stmt_2175__exit__
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237__entry__
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Update/cr
      -- 
    rr_5828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2207_inst_req_0); -- 
    cr_5833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2207_inst_req_1); -- 
    rr_5842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2211_inst_req_0); -- 
    cr_5847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2211_inst_req_1); -- 
    rr_5856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2215_inst_req_0); -- 
    cr_5861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2215_inst_req_1); -- 
    rr_5870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2219_inst_req_0); -- 
    cr_5875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(34), ack => type_cast_2219_inst_req_1); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(23) & convTransposeC_CP_5553_elements(27) & convTransposeC_CP_5553_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Sample/ra
      -- 
    ra_5829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2207_inst_ack_0, ack => convTransposeC_CP_5553_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2207_Update/ca
      -- 
    ca_5834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2207_inst_ack_1, ack => convTransposeC_CP_5553_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Sample/ra
      -- 
    ra_5843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2211_inst_ack_0, ack => convTransposeC_CP_5553_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2211_Update/ca
      -- 
    ca_5848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2211_inst_ack_1, ack => convTransposeC_CP_5553_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Sample/ra
      -- 
    ra_5857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2215_inst_ack_0, ack => convTransposeC_CP_5553_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2215_Update/ca
      -- 
    ca_5862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2215_inst_ack_1, ack => convTransposeC_CP_5553_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Sample/ra
      -- 
    ra_5871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2219_inst_ack_0, ack => convTransposeC_CP_5553_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/type_cast_2219_Update/ca
      -- 
    ca_5876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2219_inst_ack_1, ack => convTransposeC_CP_5553_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237__exit__
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2114/assign_stmt_2182_to_assign_stmt_2237/$exit
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2247/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2254/$entry
      -- CP-element group 43: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/$entry
      -- 
    rr_6268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(43), ack => type_cast_2266_inst_req_0); -- 
    cr_6273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(43), ack => type_cast_2266_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(36) & convTransposeC_CP_5553_elements(38) & convTransposeC_CP_5553_elements(40) & convTransposeC_CP_5553_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Sample/ra
      -- 
    ra_5888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2301_inst_ack_0, ack => convTransposeC_CP_5553_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Update/ca
      -- 
    ca_5893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2301_inst_ack_1, ack => convTransposeC_CP_5553_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Sample/ra
      -- 
    ra_5902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_0, ack => convTransposeC_CP_5553_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Update/ca
      -- 
    ca_5907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_1, ack => convTransposeC_CP_5553_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Sample/ra
      -- 
    ra_5916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_0, ack => convTransposeC_CP_5553_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Update/ca
      -- 
    ca_5921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_1, ack => convTransposeC_CP_5553_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Sample/ra
      -- 
    ra_5930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2339_inst_ack_0, ack => convTransposeC_CP_5553_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Sample/req
      -- 
    ca_5935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2339_inst_ack_1, ack => convTransposeC_CP_5553_elements(51)); -- 
    req_5960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(51), ack => array_obj_ref_2345_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Sample/ack
      -- 
    ack_5961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2345_index_offset_ack_0, ack => convTransposeC_CP_5553_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_request/req
      -- 
    ack_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2345_index_offset_ack_1, ack => convTransposeC_CP_5553_elements(53)); -- 
    req_5975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(53), ack => addr_of_2346_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_request/ack
      -- 
    ack_5976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2346_final_reg_ack_0, ack => convTransposeC_CP_5553_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/word_access_start/word_0/rr
      -- 
    ack_5981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2346_final_reg_ack_1, ack => convTransposeC_CP_5553_elements(55)); -- 
    rr_6014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(55), ack => ptr_deref_2350_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Sample/word_access_start/word_0/ra
      -- 
    ra_6015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2350_load_0_ack_0, ack => convTransposeC_CP_5553_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/ptr_deref_2350_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/ptr_deref_2350_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/ptr_deref_2350_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/ptr_deref_2350_Merge/merge_ack
      -- 
    ca_6026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2350_load_0_ack_1, ack => convTransposeC_CP_5553_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_index_resize_1/index_resize_ack
      -- 
    req_6056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(58), ack => array_obj_ref_2368_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(45) & convTransposeC_CP_5553_elements(47) & convTransposeC_CP_5553_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_sample_complete
      -- 
    ack_6057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2368_index_offset_ack_0, ack => convTransposeC_CP_5553_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_request/req
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_offset_calculated
      -- 
    ack_6062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2368_index_offset_ack_1, ack => convTransposeC_CP_5553_elements(60)); -- 
    req_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(60), ack => addr_of_2369_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_request/ack
      -- CP-element group 61: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_sample_completed_
      -- 
    ack_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2369_final_reg_ack_0, ack => convTransposeC_CP_5553_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_update_completed_
      -- 
    ack_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2369_final_reg_ack_1, ack => convTransposeC_CP_5553_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/ptr_deref_2372_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/ptr_deref_2372_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/ptr_deref_2372_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/ptr_deref_2372_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/$entry
      -- 
    rr_6115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(63), ack => ptr_deref_2372_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(57) & convTransposeC_CP_5553_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/word_access_start/word_0/ra
      -- CP-element group 64: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Sample/$exit
      -- 
    ra_6116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2372_store_0_ack_0, ack => convTransposeC_CP_5553_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/word_access_complete/word_0/ca
      -- 
    ca_6127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2372_store_0_ack_1, ack => convTransposeC_CP_5553_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Sample/ra
      -- 
    ra_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2377_inst_ack_0, ack => convTransposeC_CP_5553_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Update/$exit
      -- 
    ca_6141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2377_inst_ack_1, ack => convTransposeC_CP_5553_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389__exit__
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390__entry__
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2114/R_cmp_2391_place
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390_else_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2114/if_stmt_2390_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/$exit
      -- 
    branch_req_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(68), ack => if_stmt_2390_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(52) & convTransposeC_CP_5553_elements(59) & convTransposeC_CP_5553_elements(65) & convTransposeC_CP_5553_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2114/assign_stmt_2402__exit__
      -- CP-element group 69: 	 branch_block_stmt_2114/assign_stmt_2402/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2114/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2114/merge_stmt_2396__exit__
      -- CP-element group 69: 	 branch_block_stmt_2114/if_stmt_2390_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2114/assign_stmt_2402__entry__
      -- CP-element group 69: 	 branch_block_stmt_2114/assign_stmt_2402/$exit
      -- CP-element group 69: 	 branch_block_stmt_2114/if_stmt_2390_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2114/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2114/merge_stmt_2396_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2114/merge_stmt_2396_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/merge_stmt_2396_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2114/merge_stmt_2396_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2390_branch_ack_1, ack => convTransposeC_CP_5553_elements(69)); -- 
    rr_6486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(69), ack => type_cast_2454_inst_req_0); -- 
    cr_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(69), ack => type_cast_2454_inst_req_1); -- 
    rr_6509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(69), ack => type_cast_2460_inst_req_0); -- 
    cr_6514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(69), ack => type_cast_2460_inst_req_1); -- 
    rr_6532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(69), ack => type_cast_2466_inst_req_0); -- 
    cr_6537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(69), ack => type_cast_2466_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440__entry__
      -- CP-element group 70: 	 branch_block_stmt_2114/if_stmt_2390_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2114/merge_stmt_2404__exit__
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2114/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2114/if_stmt_2390_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/$entry
      -- CP-element group 70: 	 branch_block_stmt_2114/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2114/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2114/merge_stmt_2404_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2114/merge_stmt_2404_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2114/merge_stmt_2404_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2114/merge_stmt_2404_PhiAck/dummy
      -- 
    else_choice_transition_6158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2390_branch_ack_0, ack => convTransposeC_CP_5553_elements(70)); -- 
    cr_6179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(70), ack => type_cast_2418_inst_req_1); -- 
    cr_6193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(70), ack => type_cast_2434_inst_req_1); -- 
    rr_6174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(70), ack => type_cast_2418_inst_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_sample_completed_
      -- 
    ra_6175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2418_inst_ack_0, ack => convTransposeC_CP_5553_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2418_update_completed_
      -- 
    ca_6180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2418_inst_ack_1, ack => convTransposeC_CP_5553_elements(72)); -- 
    rr_6188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(72), ack => type_cast_2434_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Sample/$exit
      -- 
    ra_6189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2434_inst_ack_0, ack => convTransposeC_CP_5553_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441__entry__
      -- CP-element group 74: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440__exit__
      -- CP-element group 74: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/$exit
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2114/R_cmp122_2442_place
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2114/assign_stmt_2410_to_assign_stmt_2440/type_cast_2434_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2114/if_stmt_2441_eval_test/branch_req
      -- 
    ca_6194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2434_inst_ack_1, ack => convTransposeC_CP_5553_elements(74)); -- 
    branch_req_6202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(74), ack => if_stmt_2441_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2114/assign_stmt_2480__entry__
      -- CP-element group 75: 	 branch_block_stmt_2114/merge_stmt_2475__exit__
      -- CP-element group 75: 	 branch_block_stmt_2114/assign_stmt_2480/$entry
      -- CP-element group 75: 	 branch_block_stmt_2114/if_stmt_2441_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2114/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2114/if_stmt_2441_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2114/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2114/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2114/merge_stmt_2475_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2114/merge_stmt_2475_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2114/merge_stmt_2475_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2114/merge_stmt_2475_PhiAck/dummy
      -- 
    if_choice_transition_6207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2441_branch_ack_1, ack => convTransposeC_CP_5553_elements(75)); -- 
    req_6227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(75), ack => WPIPE_Block2_done_2477_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2114/if_stmt_2441_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2114/if_stmt_2441_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2448/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2441_branch_ack_0, ack => convTransposeC_CP_5553_elements(76)); -- 
    rr_6437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(76), ack => type_cast_2458_inst_req_0); -- 
    cr_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(76), ack => type_cast_2458_inst_req_1); -- 
    rr_6460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(76), ack => type_cast_2464_inst_req_0); -- 
    cr_6465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(76), ack => type_cast_2464_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Update/req
      -- 
    ack_6228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2477_inst_ack_0, ack => convTransposeC_CP_5553_elements(77)); -- 
    req_6232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(77), ack => WPIPE_Block2_done_2477_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2114/assign_stmt_2480__exit__
      -- CP-element group 78: 	 branch_block_stmt_2114/return__
      -- CP-element group 78: 	 branch_block_stmt_2114/merge_stmt_2482__exit__
      -- CP-element group 78: 	 branch_block_stmt_2114/branch_block_stmt_2114__exit__
      -- CP-element group 78: 	 branch_block_stmt_2114/$exit
      -- CP-element group 78: 	 branch_block_stmt_2114/assign_stmt_2480/$exit
      -- CP-element group 78: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2114/assign_stmt_2480/WPIPE_Block2_done_2477_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2114/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2114/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2114/merge_stmt_2482_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2114/merge_stmt_2482_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2114/merge_stmt_2482_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2114/merge_stmt_2482_PhiAck/dummy
      -- 
    ack_6233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2477_inst_ack_1, ack => convTransposeC_CP_5553_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 79: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2244_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- 
    phi_stmt_2240_req_6244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_6244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(79), ack => phi_stmt_2240_req_0); -- 
    -- Element group convTransposeC_CP_5553_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5553_elements(43), ack => convTransposeC_CP_5553_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2247/$exit
      -- CP-element group 80: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2251_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_req
      -- 
    phi_stmt_2247_req_6252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2247_req_6252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(80), ack => phi_stmt_2247_req_0); -- 
    -- Element group convTransposeC_CP_5553_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5553_elements(43), ack => convTransposeC_CP_5553_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Sample/ra
      -- 
    ra_6269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2266_inst_ack_0, ack => convTransposeC_CP_5553_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/Update/ca
      -- 
    ca_6274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2266_inst_ack_1, ack => convTransposeC_CP_5553_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/$exit
      -- CP-element group 83: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/$exit
      -- CP-element group 83: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2266/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_req
      -- 
    phi_stmt_2261_req_6275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2261_req_6275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(83), ack => phi_stmt_2261_req_1); -- 
    convTransposeC_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(81) & convTransposeC_CP_5553_elements(82);
      gj_convTransposeC_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2254/$exit
      -- CP-element group 84: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2258_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_req
      -- 
    phi_stmt_2254_req_6283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2254_req_6283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(84), ack => phi_stmt_2254_req_0); -- 
    -- Element group convTransposeC_CP_5553_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeC_CP_5553_elements(43), ack => convTransposeC_CP_5553_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2114/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(79) & convTransposeC_CP_5553_elements(80) & convTransposeC_CP_5553_elements(83) & convTransposeC_CP_5553_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Sample/ra
      -- 
    ra_6303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2246_inst_ack_0, ack => convTransposeC_CP_5553_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/Update/ca
      -- 
    ca_6308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2246_inst_ack_1, ack => convTransposeC_CP_5553_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 88: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/$exit
      -- CP-element group 88: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- 
    phi_stmt_2240_req_6309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_6309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(88), ack => phi_stmt_2240_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(86) & convTransposeC_CP_5553_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Sample/ra
      -- 
    ra_6326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_0, ack => convTransposeC_CP_5553_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/Update/ca
      -- 
    ca_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_1, ack => convTransposeC_CP_5553_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/$exit
      -- CP-element group 91: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/$exit
      -- CP-element group 91: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_sources/type_cast_2253/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2247/phi_stmt_2247_req
      -- 
    phi_stmt_2247_req_6332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2247_req_6332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(91), ack => phi_stmt_2247_req_1); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(89) & convTransposeC_CP_5553_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Sample/ra
      -- 
    ra_6349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2264_inst_ack_0, ack => convTransposeC_CP_5553_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/Update/ca
      -- 
    ca_6354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2264_inst_ack_1, ack => convTransposeC_CP_5553_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/$exit
      -- CP-element group 94: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/$exit
      -- CP-element group 94: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_sources/type_cast_2264/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2261/phi_stmt_2261_req
      -- 
    phi_stmt_2261_req_6355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2261_req_6355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(94), ack => phi_stmt_2261_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(92) & convTransposeC_CP_5553_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Sample/ra
      -- 
    ra_6372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_0, ack => convTransposeC_CP_5553_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/Update/ca
      -- 
    ca_6377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_1, ack => convTransposeC_CP_5553_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/$exit
      -- CP-element group 97: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/$exit
      -- CP-element group 97: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_sources/type_cast_2260/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2254/phi_stmt_2254_req
      -- 
    phi_stmt_2254_req_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2254_req_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(97), ack => phi_stmt_2254_req_1); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(95) & convTransposeC_CP_5553_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2114/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(88) & convTransposeC_CP_5553_elements(91) & convTransposeC_CP_5553_elements(94) & convTransposeC_CP_5553_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2114/merge_stmt_2239_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2114/merge_stmt_2239_PhiAck/$entry
      -- 
    convTransposeC_CP_5553_elements(99) <= OrReduce(convTransposeC_CP_5553_elements(85) & convTransposeC_CP_5553_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2114/merge_stmt_2239_PhiAck/phi_stmt_2240_ack
      -- 
    phi_stmt_2240_ack_6383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2240_ack_0, ack => convTransposeC_CP_5553_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2114/merge_stmt_2239_PhiAck/phi_stmt_2247_ack
      -- 
    phi_stmt_2247_ack_6384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2247_ack_0, ack => convTransposeC_CP_5553_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2114/merge_stmt_2239_PhiAck/phi_stmt_2254_ack
      -- 
    phi_stmt_2254_ack_6385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2254_ack_0, ack => convTransposeC_CP_5553_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2114/merge_stmt_2239_PhiAck/phi_stmt_2261_ack
      -- 
    phi_stmt_2261_ack_6386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2261_ack_0, ack => convTransposeC_CP_5553_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/merge_stmt_2239__exit__
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389__entry__
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2372_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2368_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2377_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2301_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2305_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2309_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/type_cast_2339_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/array_obj_ref_2345_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2346_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/ptr_deref_2350_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2114/assign_stmt_2273_to_assign_stmt_2389/addr_of_2369_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2114/merge_stmt_2239_PhiAck/$exit
      -- 
    req_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => addr_of_2369_final_reg_req_1); -- 
    cr_6126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => ptr_deref_2372_store_0_req_1); -- 
    rr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2377_inst_req_0); -- 
    req_6061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => array_obj_ref_2368_index_offset_req_1); -- 
    cr_6140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2377_inst_req_1); -- 
    rr_5887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2301_inst_req_0); -- 
    cr_5892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2301_inst_req_1); -- 
    rr_5901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2305_inst_req_0); -- 
    cr_5906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2305_inst_req_1); -- 
    rr_5915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2309_inst_req_0); -- 
    cr_5920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2309_inst_req_1); -- 
    rr_5929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2339_inst_req_0); -- 
    cr_5934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => type_cast_2339_inst_req_1); -- 
    req_5965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => array_obj_ref_2345_index_offset_req_1); -- 
    req_5980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => addr_of_2346_final_reg_req_1); -- 
    cr_6025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(104), ack => ptr_deref_2350_load_0_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(100) & convTransposeC_CP_5553_elements(101) & convTransposeC_CP_5553_elements(102) & convTransposeC_CP_5553_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2448/$exit
      -- CP-element group 105: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2452_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_req
      -- 
    phi_stmt_2448_req_6421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2448_req_6421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(105), ack => phi_stmt_2448_req_0); -- 
    -- Element group convTransposeC_CP_5553_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5553_elements(76), ack => convTransposeC_CP_5553_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Sample/ra
      -- 
    ra_6438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2458_inst_ack_0, ack => convTransposeC_CP_5553_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/Update/ca
      -- 
    ca_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2458_inst_ack_1, ack => convTransposeC_CP_5553_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/$exit
      -- CP-element group 108: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/$exit
      -- CP-element group 108: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2458/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_req
      -- 
    phi_stmt_2455_req_6444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2455_req_6444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(108), ack => phi_stmt_2455_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(106) & convTransposeC_CP_5553_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Sample/ra
      -- 
    ra_6461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2464_inst_ack_0, ack => convTransposeC_CP_5553_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/Update/ca
      -- 
    ca_6466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2464_inst_ack_1, ack => convTransposeC_CP_5553_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/$exit
      -- CP-element group 111: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/$exit
      -- CP-element group 111: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2464/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_req
      -- 
    phi_stmt_2461_req_6467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2461_req_6467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(111), ack => phi_stmt_2461_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(109) & convTransposeC_CP_5553_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2114/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(105) & convTransposeC_CP_5553_elements(108) & convTransposeC_CP_5553_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Sample/ra
      -- 
    ra_6487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2454_inst_ack_0, ack => convTransposeC_CP_5553_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/Update/ca
      -- 
    ca_6492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2454_inst_ack_1, ack => convTransposeC_CP_5553_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/$exit
      -- CP-element group 115: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/$exit
      -- CP-element group 115: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_sources/type_cast_2454/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2448/phi_stmt_2448_req
      -- 
    phi_stmt_2448_req_6493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2448_req_6493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(115), ack => phi_stmt_2448_req_1); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(113) & convTransposeC_CP_5553_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Sample/ra
      -- 
    ra_6510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_0, ack => convTransposeC_CP_5553_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/Update/ca
      -- 
    ca_6515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_1, ack => convTransposeC_CP_5553_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/$exit
      -- CP-element group 118: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/$exit
      -- CP-element group 118: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_sources/type_cast_2460/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2455/phi_stmt_2455_req
      -- 
    phi_stmt_2455_req_6516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2455_req_6516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(118), ack => phi_stmt_2455_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(116) & convTransposeC_CP_5553_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Sample/ra
      -- 
    ra_6533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2466_inst_ack_0, ack => convTransposeC_CP_5553_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/Update/ca
      -- 
    ca_6538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2466_inst_ack_1, ack => convTransposeC_CP_5553_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/$exit
      -- CP-element group 121: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/$exit
      -- CP-element group 121: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_sources/type_cast_2466/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2461/phi_stmt_2461_req
      -- 
    phi_stmt_2461_req_6539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2461_req_6539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5553_elements(121), ack => phi_stmt_2461_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(119) & convTransposeC_CP_5553_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2114/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(115) & convTransposeC_CP_5553_elements(118) & convTransposeC_CP_5553_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2114/merge_stmt_2447_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2114/merge_stmt_2447_PhiAck/$entry
      -- 
    convTransposeC_CP_5553_elements(123) <= OrReduce(convTransposeC_CP_5553_elements(112) & convTransposeC_CP_5553_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2114/merge_stmt_2447_PhiAck/phi_stmt_2448_ack
      -- 
    phi_stmt_2448_ack_6544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2448_ack_0, ack => convTransposeC_CP_5553_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2114/merge_stmt_2447_PhiAck/phi_stmt_2455_ack
      -- 
    phi_stmt_2455_ack_6545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2455_ack_0, ack => convTransposeC_CP_5553_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2114/merge_stmt_2447_PhiAck/phi_stmt_2461_ack
      -- 
    phi_stmt_2461_ack_6546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2461_ack_0, ack => convTransposeC_CP_5553_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2114/merge_stmt_2447_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5553_elements(124) & convTransposeC_CP_5553_elements(125) & convTransposeC_CP_5553_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5553_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2367_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2367_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2344_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2344_scaled : std_logic_vector(13 downto 0);
    signal add121_2237 : std_logic_vector(31 downto 0);
    signal add45_2188 : std_logic_vector(15 downto 0);
    signal add58_2199 : std_logic_vector(15 downto 0);
    signal add77_2320 : std_logic_vector(63 downto 0);
    signal add79_2330 : std_logic_vector(63 downto 0);
    signal add91_2384 : std_logic_vector(31 downto 0);
    signal add98_2402 : std_logic_vector(15 downto 0);
    signal add_2166 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2278 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2345_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2345_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2345_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2345_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2345_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2345_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2368_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2368_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2368_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2368_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2368_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2368_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2347 : std_logic_vector(31 downto 0);
    signal arrayidx87_2370 : std_logic_vector(31 downto 0);
    signal call11_2135 : std_logic_vector(15 downto 0);
    signal call13_2138 : std_logic_vector(15 downto 0);
    signal call14_2141 : std_logic_vector(15 downto 0);
    signal call15_2144 : std_logic_vector(15 downto 0);
    signal call16_2157 : std_logic_vector(15 downto 0);
    signal call18_2169 : std_logic_vector(15 downto 0);
    signal call1_2120 : std_logic_vector(15 downto 0);
    signal call20_2172 : std_logic_vector(15 downto 0);
    signal call22_2175 : std_logic_vector(15 downto 0);
    signal call3_2123 : std_logic_vector(15 downto 0);
    signal call5_2126 : std_logic_vector(15 downto 0);
    signal call7_2129 : std_logic_vector(15 downto 0);
    signal call9_2132 : std_logic_vector(15 downto 0);
    signal call_2117 : std_logic_vector(15 downto 0);
    signal cmp106_2415 : std_logic_vector(0 downto 0);
    signal cmp122_2440 : std_logic_vector(0 downto 0);
    signal cmp_2389 : std_logic_vector(0 downto 0);
    signal conv112_2435 : std_logic_vector(31 downto 0);
    signal conv115_2220 : std_logic_vector(31 downto 0);
    signal conv17_2161 : std_logic_vector(31 downto 0);
    signal conv65_2302 : std_logic_vector(63 downto 0);
    signal conv68_2208 : std_logic_vector(63 downto 0);
    signal conv70_2306 : std_logic_vector(63 downto 0);
    signal conv73_2212 : std_logic_vector(63 downto 0);
    signal conv75_2310 : std_logic_vector(63 downto 0);
    signal conv90_2378 : std_logic_vector(31 downto 0);
    signal conv94_2216 : std_logic_vector(31 downto 0);
    signal conv_2148 : std_logic_vector(31 downto 0);
    signal idxprom86_2363 : std_logic_vector(63 downto 0);
    signal idxprom_2340 : std_logic_vector(63 downto 0);
    signal inc110_2419 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2424 : std_logic_vector(15 downto 0);
    signal inc_2410 : std_logic_vector(15 downto 0);
    signal indvar_2240 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2473 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2461 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2261 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2455 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2254 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2431 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2448 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2247 : std_logic_vector(15 downto 0);
    signal mul54_2293 : std_logic_vector(15 downto 0);
    signal mul76_2315 : std_logic_vector(63 downto 0);
    signal mul78_2325 : std_logic_vector(63 downto 0);
    signal mul_2283 : std_logic_vector(15 downto 0);
    signal ptr_deref_2350_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2350_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2350_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2350_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2350_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2372_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2372_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2372_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2372_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2372_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2372_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2154 : std_logic_vector(31 downto 0);
    signal shr116137_2226 : std_logic_vector(31 downto 0);
    signal shr120138_2232 : std_logic_vector(31 downto 0);
    signal shr136_2182 : std_logic_vector(15 downto 0);
    signal shr81_2336 : std_logic_vector(31 downto 0);
    signal shr85_2357 : std_logic_vector(63 downto 0);
    signal sub48_2288 : std_logic_vector(15 downto 0);
    signal sub61_2204 : std_logic_vector(15 downto 0);
    signal sub62_2298 : std_logic_vector(15 downto 0);
    signal sub_2193 : std_logic_vector(15 downto 0);
    signal tmp1_2273 : std_logic_vector(31 downto 0);
    signal tmp83_2351 : std_logic_vector(63 downto 0);
    signal type_cast_2152_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2180_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2186_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2197_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2224_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2230_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2244_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2246_wire : std_logic_vector(31 downto 0);
    signal type_cast_2251_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2253_wire : std_logic_vector(15 downto 0);
    signal type_cast_2258_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2260_wire : std_logic_vector(15 downto 0);
    signal type_cast_2264_wire : std_logic_vector(15 downto 0);
    signal type_cast_2266_wire : std_logic_vector(15 downto 0);
    signal type_cast_2271_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2334_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2355_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2361_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2382_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2400_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2408_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2428_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2452_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2454_wire : std_logic_vector(15 downto 0);
    signal type_cast_2458_wire : std_logic_vector(15 downto 0);
    signal type_cast_2460_wire : std_logic_vector(15 downto 0);
    signal type_cast_2464_wire : std_logic_vector(15 downto 0);
    signal type_cast_2466_wire : std_logic_vector(15 downto 0);
    signal type_cast_2471_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2479_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2345_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2345_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2345_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2345_resized_base_address <= "00000000000000";
    array_obj_ref_2368_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2368_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2368_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2368_resized_base_address <= "00000000000000";
    ptr_deref_2350_word_offset_0 <= "00000000000000";
    ptr_deref_2372_word_offset_0 <= "00000000000000";
    type_cast_2152_wire_constant <= "00000000000000000000000000010000";
    type_cast_2180_wire_constant <= "0000000000000001";
    type_cast_2186_wire_constant <= "1111111111111111";
    type_cast_2197_wire_constant <= "1111111111111111";
    type_cast_2224_wire_constant <= "00000000000000000000000000000010";
    type_cast_2230_wire_constant <= "00000000000000000000000000000001";
    type_cast_2244_wire_constant <= "00000000000000000000000000000000";
    type_cast_2251_wire_constant <= "0000000000000000";
    type_cast_2258_wire_constant <= "0000000000000000";
    type_cast_2271_wire_constant <= "00000000000000000000000000000100";
    type_cast_2334_wire_constant <= "00000000000000000000000000000010";
    type_cast_2355_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2361_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2382_wire_constant <= "00000000000000000000000000000100";
    type_cast_2400_wire_constant <= "0000000000000100";
    type_cast_2408_wire_constant <= "0000000000000001";
    type_cast_2428_wire_constant <= "0000000000000000";
    type_cast_2452_wire_constant <= "0000000000000000";
    type_cast_2471_wire_constant <= "00000000000000000000000000000001";
    type_cast_2479_wire_constant <= "0000000000000001";
    phi_stmt_2240: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2244_wire_constant & type_cast_2246_wire;
      req <= phi_stmt_2240_req_0 & phi_stmt_2240_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2240",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2240_ack_0,
          idata => idata,
          odata => indvar_2240,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2240
    phi_stmt_2247: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2251_wire_constant & type_cast_2253_wire;
      req <= phi_stmt_2247_req_0 & phi_stmt_2247_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2247",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2247_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2247,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2247
    phi_stmt_2254: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2258_wire_constant & type_cast_2260_wire;
      req <= phi_stmt_2254_req_0 & phi_stmt_2254_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2254",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2254_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2254,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2254
    phi_stmt_2261: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2264_wire & type_cast_2266_wire;
      req <= phi_stmt_2261_req_0 & phi_stmt_2261_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2261",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2261_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2261,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2261
    phi_stmt_2448: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2452_wire_constant & type_cast_2454_wire;
      req <= phi_stmt_2448_req_0 & phi_stmt_2448_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2448",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2448_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2448,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2448
    phi_stmt_2455: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2458_wire & type_cast_2460_wire;
      req <= phi_stmt_2455_req_0 & phi_stmt_2455_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2455",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2455_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2455,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2455
    phi_stmt_2461: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2464_wire & type_cast_2466_wire;
      req <= phi_stmt_2461_req_0 & phi_stmt_2461_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2461",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2461_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2461,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2461
    -- flow-through select operator MUX_2430_inst
    input_dim1x_x2_2431 <= type_cast_2428_wire_constant when (cmp106_2415(0) /=  '0') else inc_2410;
    addr_of_2346_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2346_final_reg_req_0;
      addr_of_2346_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2346_final_reg_req_1;
      addr_of_2346_final_reg_ack_1<= rack(0);
      addr_of_2346_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2346_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2345_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2369_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2369_final_reg_req_0;
      addr_of_2369_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2369_final_reg_req_1;
      addr_of_2369_final_reg_ack_1<= rack(0);
      addr_of_2369_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2369_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2368_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2147_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2147_inst_req_0;
      type_cast_2147_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2147_inst_req_1;
      type_cast_2147_inst_ack_1<= rack(0);
      type_cast_2147_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2147_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2148,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2160_inst_req_0;
      type_cast_2160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2160_inst_req_1;
      type_cast_2160_inst_ack_1<= rack(0);
      type_cast_2160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2207_inst_req_0;
      type_cast_2207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2207_inst_req_1;
      type_cast_2207_inst_ack_1<= rack(0);
      type_cast_2207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2211_inst_req_0;
      type_cast_2211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2211_inst_req_1;
      type_cast_2211_inst_ack_1<= rack(0);
      type_cast_2211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2172,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2215_inst_req_0;
      type_cast_2215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2215_inst_req_1;
      type_cast_2215_inst_ack_1<= rack(0);
      type_cast_2215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2219_inst_req_0;
      type_cast_2219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2219_inst_req_1;
      type_cast_2219_inst_ack_1<= rack(0);
      type_cast_2219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2246_inst_req_0;
      type_cast_2246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2246_inst_req_1;
      type_cast_2246_inst_ack_1<= rack(0);
      type_cast_2246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2473,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2246_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2253_inst_req_0;
      type_cast_2253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2253_inst_req_1;
      type_cast_2253_inst_ack_1<= rack(0);
      type_cast_2253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2253_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2260_inst_req_0;
      type_cast_2260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2260_inst_req_1;
      type_cast_2260_inst_ack_1<= rack(0);
      type_cast_2260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2260_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2264_inst_req_0;
      type_cast_2264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2264_inst_req_1;
      type_cast_2264_inst_ack_1<= rack(0);
      type_cast_2264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2461,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2264_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2266_inst_req_0;
      type_cast_2266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2266_inst_req_1;
      type_cast_2266_inst_ack_1<= rack(0);
      type_cast_2266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2266_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2301_inst_req_0;
      type_cast_2301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2301_inst_req_1;
      type_cast_2301_inst_ack_1<= rack(0);
      type_cast_2301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2305_inst_req_0;
      type_cast_2305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2305_inst_req_1;
      type_cast_2305_inst_ack_1<= rack(0);
      type_cast_2305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2309_inst_req_0;
      type_cast_2309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2309_inst_req_1;
      type_cast_2309_inst_ack_1<= rack(0);
      type_cast_2309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2339_inst_req_0;
      type_cast_2339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2339_inst_req_1;
      type_cast_2339_inst_ack_1<= rack(0);
      type_cast_2339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2377_inst_req_0;
      type_cast_2377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2377_inst_req_1;
      type_cast_2377_inst_ack_1<= rack(0);
      type_cast_2377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2418_inst_req_0;
      type_cast_2418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2418_inst_req_1;
      type_cast_2418_inst_ack_1<= rack(0);
      type_cast_2418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2434_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2434_inst_req_0;
      type_cast_2434_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2434_inst_req_1;
      type_cast_2434_inst_ack_1<= rack(0);
      type_cast_2434_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2434_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2435,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2454_inst_req_0;
      type_cast_2454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2454_inst_req_1;
      type_cast_2454_inst_ack_1<= rack(0);
      type_cast_2454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2454_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2458_inst_req_0;
      type_cast_2458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2458_inst_req_1;
      type_cast_2458_inst_ack_1<= rack(0);
      type_cast_2458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2431,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2458_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2460_inst_req_0;
      type_cast_2460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2460_inst_req_1;
      type_cast_2460_inst_ack_1<= rack(0);
      type_cast_2460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2460_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2464_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2464_inst_req_0;
      type_cast_2464_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2464_inst_req_1;
      type_cast_2464_inst_ack_1<= rack(0);
      type_cast_2464_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2464_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2464_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2466_inst_req_0;
      type_cast_2466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2466_inst_req_1;
      type_cast_2466_inst_ack_1<= rack(0);
      type_cast_2466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2261,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2466_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2345_index_1_rename
    process(R_idxprom_2344_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2344_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2344_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2345_index_1_resize
    process(idxprom_2340) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2340;
      ov := iv(13 downto 0);
      R_idxprom_2344_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2345_root_address_inst
    process(array_obj_ref_2345_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2345_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2345_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2368_index_1_rename
    process(R_idxprom86_2367_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2367_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2367_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2368_index_1_resize
    process(idxprom86_2363) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2363;
      ov := iv(13 downto 0);
      R_idxprom86_2367_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2368_root_address_inst
    process(array_obj_ref_2368_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2368_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2368_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_addr_0
    process(ptr_deref_2350_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2350_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2350_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_base_resize
    process(arrayidx82_2347) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2347;
      ov := iv(13 downto 0);
      ptr_deref_2350_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_gather_scatter
    process(ptr_deref_2350_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2350_data_0;
      ov(63 downto 0) := iv;
      tmp83_2351 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2350_root_address_inst
    process(ptr_deref_2350_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2350_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2350_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_addr_0
    process(ptr_deref_2372_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2372_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2372_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_base_resize
    process(arrayidx87_2370) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2370;
      ov := iv(13 downto 0);
      ptr_deref_2372_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_gather_scatter
    process(tmp83_2351) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2351;
      ov(63 downto 0) := iv;
      ptr_deref_2372_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2372_root_address_inst
    process(ptr_deref_2372_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2372_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2372_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2390_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2389;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2390_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2390_branch_req_0,
          ack0 => if_stmt_2390_branch_ack_0,
          ack1 => if_stmt_2390_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2441_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2440;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2441_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2441_branch_req_0,
          ack0 => if_stmt_2441_branch_ack_0,
          ack1 => if_stmt_2441_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2187_inst
    process(call7_2129) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2129, type_cast_2186_wire_constant, tmp_var);
      add45_2188 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2198_inst
    process(call9_2132) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2132, type_cast_2197_wire_constant, tmp_var);
      add58_2199 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2287_inst
    process(sub_2193, mul_2283) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2193, mul_2283, tmp_var);
      sub48_2288 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2297_inst
    process(sub61_2204, mul54_2293) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2204, mul54_2293, tmp_var);
      sub62_2298 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2401_inst
    process(input_dim2x_x1_2247) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2247, type_cast_2400_wire_constant, tmp_var);
      add98_2402 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2409_inst
    process(input_dim1x_x1_2254) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2254, type_cast_2408_wire_constant, tmp_var);
      inc_2410 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2423_inst
    process(inc110_2419, input_dim0x_x2_2261) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2419, input_dim0x_x2_2261, tmp_var);
      inc110x_xinput_dim0x_x2_2424 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2236_inst
    process(shr116137_2226, shr120138_2232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2226, shr120138_2232, tmp_var);
      add121_2237 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2277_inst
    process(add_2166, tmp1_2273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2166, tmp1_2273, tmp_var);
      add_src_0x_x0_2278 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2383_inst
    process(conv90_2378) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2378, type_cast_2382_wire_constant, tmp_var);
      add91_2384 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2472_inst
    process(indvar_2240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2240, type_cast_2471_wire_constant, tmp_var);
      indvarx_xnext_2473 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2319_inst
    process(mul76_2315, conv70_2306) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2315, conv70_2306, tmp_var);
      add77_2320 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2329_inst
    process(mul78_2325, conv65_2302) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2325, conv65_2302, tmp_var);
      add79_2330 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2362_inst
    process(shr85_2357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2357, type_cast_2361_wire_constant, tmp_var);
      idxprom86_2363 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2414_inst
    process(inc_2410, call1_2120) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2410, call1_2120, tmp_var);
      cmp106_2415 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2439_inst
    process(conv112_2435, add121_2237) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2435, add121_2237, tmp_var);
      cmp122_2440 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2181_inst
    process(call_2117) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2117, type_cast_2180_wire_constant, tmp_var);
      shr136_2182 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2225_inst
    process(conv115_2220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2220, type_cast_2224_wire_constant, tmp_var);
      shr116137_2226 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2231_inst
    process(conv115_2220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2220, type_cast_2230_wire_constant, tmp_var);
      shr120138_2232 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2335_inst
    process(add_src_0x_x0_2278) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2278, type_cast_2334_wire_constant, tmp_var);
      shr81_2336 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2356_inst
    process(add79_2330) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2330, type_cast_2355_wire_constant, tmp_var);
      shr85_2357 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2282_inst
    process(input_dim0x_x2_2261, call13_2138) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2261, call13_2138, tmp_var);
      mul_2283 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2292_inst
    process(input_dim1x_x1_2254, call13_2138) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2254, call13_2138, tmp_var);
      mul54_2293 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2272_inst
    process(indvar_2240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2240, type_cast_2271_wire_constant, tmp_var);
      tmp1_2273 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2314_inst
    process(conv75_2310, conv73_2212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2310, conv73_2212, tmp_var);
      mul76_2315 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2324_inst
    process(add77_2320, conv68_2208) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2320, conv68_2208, tmp_var);
      mul78_2325 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2165_inst
    process(shl_2154, conv17_2161) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2154, conv17_2161, tmp_var);
      add_2166 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2153_inst
    process(conv_2148) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2148, type_cast_2152_wire_constant, tmp_var);
      shl_2154 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2192_inst
    process(add45_2188, call14_2141) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2188, call14_2141, tmp_var);
      sub_2193 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2203_inst
    process(add58_2199, call14_2141) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2199, call14_2141, tmp_var);
      sub61_2204 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2388_inst
    process(add91_2384, conv94_2216) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2384, conv94_2216, tmp_var);
      cmp_2389 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2345_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2344_scaled;
      array_obj_ref_2345_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2345_index_offset_req_0;
      array_obj_ref_2345_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2345_index_offset_req_1;
      array_obj_ref_2345_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2368_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2367_scaled;
      array_obj_ref_2368_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2368_index_offset_req_0;
      array_obj_ref_2368_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2368_index_offset_req_1;
      array_obj_ref_2368_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2350_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2350_load_0_req_0;
      ptr_deref_2350_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2350_load_0_req_1;
      ptr_deref_2350_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2350_word_address_0;
      ptr_deref_2350_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2372_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2372_store_0_req_0;
      ptr_deref_2372_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2372_store_0_req_1;
      ptr_deref_2372_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2372_word_address_0;
      data_in <= ptr_deref_2372_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2116_inst RPIPE_Block2_start_2119_inst RPIPE_Block2_start_2122_inst RPIPE_Block2_start_2125_inst RPIPE_Block2_start_2128_inst RPIPE_Block2_start_2131_inst RPIPE_Block2_start_2134_inst RPIPE_Block2_start_2137_inst RPIPE_Block2_start_2140_inst RPIPE_Block2_start_2143_inst RPIPE_Block2_start_2156_inst RPIPE_Block2_start_2168_inst RPIPE_Block2_start_2171_inst RPIPE_Block2_start_2174_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2116_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2119_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2122_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2125_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2128_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2131_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2134_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2137_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2140_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2143_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2156_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2168_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2171_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2174_inst_req_0;
      RPIPE_Block2_start_2116_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2119_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2122_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2125_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2128_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2131_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2134_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2137_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2140_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2143_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2156_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2168_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2171_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2174_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2116_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2119_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2122_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2125_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2128_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2131_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2134_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2137_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2140_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2143_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2156_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2168_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2171_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2174_inst_req_1;
      RPIPE_Block2_start_2116_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2119_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2122_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2125_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2128_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2131_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2134_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2137_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2140_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2143_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2156_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2168_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2171_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2174_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2117 <= data_out(223 downto 208);
      call1_2120 <= data_out(207 downto 192);
      call3_2123 <= data_out(191 downto 176);
      call5_2126 <= data_out(175 downto 160);
      call7_2129 <= data_out(159 downto 144);
      call9_2132 <= data_out(143 downto 128);
      call11_2135 <= data_out(127 downto 112);
      call13_2138 <= data_out(111 downto 96);
      call14_2141 <= data_out(95 downto 80);
      call15_2144 <= data_out(79 downto 64);
      call16_2157 <= data_out(63 downto 48);
      call18_2169 <= data_out(47 downto 32);
      call20_2172 <= data_out(31 downto 16);
      call22_2175 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2477_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2477_inst_req_0;
      WPIPE_Block2_done_2477_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2477_inst_req_1;
      WPIPE_Block2_done_2477_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2479_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6563_start: Boolean;
  signal convTransposeD_CP_6563_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2497_inst_ack_0 : boolean;
  signal addr_of_2731_final_reg_req_0 : boolean;
  signal RPIPE_Block3_start_2503_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2503_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2491_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2500_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2491_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2503_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2491_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2491_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2503_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2497_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2497_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2494_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2494_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2488_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2488_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2494_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2494_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2488_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2488_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2500_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2500_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2500_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2497_inst_req_0 : boolean;
  signal type_cast_2615_inst_ack_1 : boolean;
  signal addr_of_2731_final_reg_ack_0 : boolean;
  signal if_stmt_2799_branch_ack_0 : boolean;
  signal type_cast_2622_inst_req_1 : boolean;
  signal type_cast_2622_inst_ack_1 : boolean;
  signal phi_stmt_2623_req_0 : boolean;
  signal phi_stmt_2609_req_1 : boolean;
  signal type_cast_2622_inst_req_0 : boolean;
  signal type_cast_2608_inst_req_0 : boolean;
  signal type_cast_2608_inst_ack_0 : boolean;
  signal type_cast_2615_inst_req_0 : boolean;
  signal type_cast_2622_inst_ack_0 : boolean;
  signal phi_stmt_2616_req_1 : boolean;
  signal type_cast_2615_inst_ack_0 : boolean;
  signal addr_of_2731_final_reg_req_1 : boolean;
  signal type_cast_2628_inst_req_0 : boolean;
  signal type_cast_2628_inst_ack_0 : boolean;
  signal addr_of_2731_final_reg_ack_1 : boolean;
  signal type_cast_2626_inst_req_0 : boolean;
  signal ptr_deref_2734_store_0_req_0 : boolean;
  signal ptr_deref_2734_store_0_ack_0 : boolean;
  signal type_cast_2628_inst_req_1 : boolean;
  signal type_cast_2628_inst_ack_1 : boolean;
  signal type_cast_2608_inst_req_1 : boolean;
  signal type_cast_2608_inst_ack_1 : boolean;
  signal phi_stmt_2616_req_0 : boolean;
  signal phi_stmt_2602_req_1 : boolean;
  signal type_cast_2626_inst_ack_0 : boolean;
  signal if_stmt_2799_branch_req_0 : boolean;
  signal if_stmt_2752_branch_ack_0 : boolean;
  signal type_cast_2780_inst_req_1 : boolean;
  signal type_cast_2626_inst_req_1 : boolean;
  signal ptr_deref_2734_store_0_req_1 : boolean;
  signal ptr_deref_2734_store_0_ack_1 : boolean;
  signal type_cast_2780_inst_ack_1 : boolean;
  signal array_obj_ref_2730_index_offset_req_0 : boolean;
  signal phi_stmt_2623_req_1 : boolean;
  signal type_cast_2615_inst_req_1 : boolean;
  signal phi_stmt_2602_ack_0 : boolean;
  signal RPIPE_Block3_start_2506_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2506_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2506_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2506_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2509_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2509_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2509_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2509_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2512_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2512_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2512_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2512_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2515_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2515_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2515_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2515_inst_ack_1 : boolean;
  signal type_cast_2519_inst_req_0 : boolean;
  signal type_cast_2519_inst_ack_0 : boolean;
  signal type_cast_2519_inst_req_1 : boolean;
  signal type_cast_2519_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2528_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2528_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2528_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2528_inst_ack_1 : boolean;
  signal type_cast_2532_inst_req_0 : boolean;
  signal type_cast_2532_inst_ack_0 : boolean;
  signal type_cast_2532_inst_req_1 : boolean;
  signal type_cast_2532_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2540_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2540_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2540_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2540_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2543_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2543_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2543_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2543_inst_ack_1 : boolean;
  signal phi_stmt_2609_req_0 : boolean;
  signal type_cast_2780_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2546_inst_req_0 : boolean;
  signal if_stmt_2752_branch_ack_1 : boolean;
  signal RPIPE_Block3_start_2546_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2546_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2546_inst_ack_1 : boolean;
  signal if_stmt_2799_branch_ack_1 : boolean;
  signal type_cast_2780_inst_req_0 : boolean;
  signal type_cast_2590_inst_req_0 : boolean;
  signal type_cast_2590_inst_ack_0 : boolean;
  signal type_cast_2590_inst_req_1 : boolean;
  signal if_stmt_2752_branch_req_0 : boolean;
  signal type_cast_2590_inst_ack_1 : boolean;
  signal type_cast_2626_inst_ack_1 : boolean;
  signal type_cast_2594_inst_req_0 : boolean;
  signal type_cast_2594_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2835_inst_ack_1 : boolean;
  signal type_cast_2594_inst_req_1 : boolean;
  signal type_cast_2594_inst_ack_1 : boolean;
  signal WPIPE_Block3_done_2835_inst_req_1 : boolean;
  signal type_cast_2598_inst_req_0 : boolean;
  signal type_cast_2598_inst_ack_0 : boolean;
  signal type_cast_2598_inst_req_1 : boolean;
  signal type_cast_2598_inst_ack_1 : boolean;
  signal phi_stmt_2602_req_0 : boolean;
  signal type_cast_2663_inst_req_0 : boolean;
  signal type_cast_2739_inst_ack_1 : boolean;
  signal type_cast_2663_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2835_inst_ack_0 : boolean;
  signal type_cast_2663_inst_req_1 : boolean;
  signal type_cast_2739_inst_req_1 : boolean;
  signal type_cast_2663_inst_ack_1 : boolean;
  signal array_obj_ref_2730_index_offset_ack_1 : boolean;
  signal WPIPE_Block3_done_2835_inst_req_0 : boolean;
  signal type_cast_2667_inst_req_0 : boolean;
  signal type_cast_2667_inst_ack_0 : boolean;
  signal type_cast_2667_inst_req_1 : boolean;
  signal type_cast_2667_inst_ack_1 : boolean;
  signal array_obj_ref_2730_index_offset_req_1 : boolean;
  signal type_cast_2671_inst_req_0 : boolean;
  signal type_cast_2739_inst_ack_0 : boolean;
  signal type_cast_2671_inst_ack_0 : boolean;
  signal type_cast_2671_inst_req_1 : boolean;
  signal type_cast_2739_inst_req_0 : boolean;
  signal type_cast_2671_inst_ack_1 : boolean;
  signal array_obj_ref_2730_index_offset_ack_0 : boolean;
  signal type_cast_2701_inst_req_0 : boolean;
  signal type_cast_2701_inst_ack_0 : boolean;
  signal type_cast_2701_inst_req_1 : boolean;
  signal type_cast_2701_inst_ack_1 : boolean;
  signal array_obj_ref_2707_index_offset_req_0 : boolean;
  signal array_obj_ref_2707_index_offset_ack_0 : boolean;
  signal array_obj_ref_2707_index_offset_req_1 : boolean;
  signal array_obj_ref_2707_index_offset_ack_1 : boolean;
  signal addr_of_2708_final_reg_req_0 : boolean;
  signal addr_of_2708_final_reg_ack_0 : boolean;
  signal addr_of_2708_final_reg_req_1 : boolean;
  signal addr_of_2708_final_reg_ack_1 : boolean;
  signal ptr_deref_2712_load_0_req_0 : boolean;
  signal ptr_deref_2712_load_0_ack_0 : boolean;
  signal ptr_deref_2712_load_0_req_1 : boolean;
  signal ptr_deref_2712_load_0_ack_1 : boolean;
  signal phi_stmt_2609_ack_0 : boolean;
  signal phi_stmt_2616_ack_0 : boolean;
  signal phi_stmt_2623_ack_0 : boolean;
  signal phi_stmt_2806_req_1 : boolean;
  signal type_cast_2818_inst_req_0 : boolean;
  signal type_cast_2818_inst_ack_0 : boolean;
  signal type_cast_2818_inst_req_1 : boolean;
  signal type_cast_2818_inst_ack_1 : boolean;
  signal phi_stmt_2813_req_1 : boolean;
  signal type_cast_2824_inst_req_0 : boolean;
  signal type_cast_2824_inst_ack_0 : boolean;
  signal type_cast_2824_inst_req_1 : boolean;
  signal type_cast_2824_inst_ack_1 : boolean;
  signal phi_stmt_2819_req_1 : boolean;
  signal type_cast_2809_inst_req_0 : boolean;
  signal type_cast_2809_inst_ack_0 : boolean;
  signal type_cast_2809_inst_req_1 : boolean;
  signal type_cast_2809_inst_ack_1 : boolean;
  signal phi_stmt_2806_req_0 : boolean;
  signal type_cast_2816_inst_req_0 : boolean;
  signal type_cast_2816_inst_ack_0 : boolean;
  signal type_cast_2816_inst_req_1 : boolean;
  signal type_cast_2816_inst_ack_1 : boolean;
  signal phi_stmt_2813_req_0 : boolean;
  signal type_cast_2822_inst_req_0 : boolean;
  signal type_cast_2822_inst_ack_0 : boolean;
  signal type_cast_2822_inst_req_1 : boolean;
  signal type_cast_2822_inst_ack_1 : boolean;
  signal phi_stmt_2819_req_0 : boolean;
  signal phi_stmt_2806_ack_0 : boolean;
  signal phi_stmt_2813_ack_0 : boolean;
  signal phi_stmt_2819_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6563_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6563_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6563_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6563_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6563: Block -- control-path 
    signal convTransposeD_CP_6563_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6563_elements(0) <= convTransposeD_CP_6563_start;
    convTransposeD_CP_6563_symbol <= convTransposeD_CP_6563_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2486/$entry
      -- CP-element group 0: 	 branch_block_stmt_2486/branch_block_stmt_2486__entry__
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547__entry__
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/$entry
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Update/cr
      -- 
    rr_6611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(0), ack => RPIPE_Block3_start_2488_inst_req_0); -- 
    cr_6756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(0), ack => type_cast_2519_inst_req_1); -- 
    cr_6784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(0), ack => type_cast_2532_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/assign_stmt_2831/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2486/assign_stmt_2831/$exit
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2486/merge_stmt_2805__exit__
      -- CP-element group 1: 	 branch_block_stmt_2486/assign_stmt_2831__entry__
      -- CP-element group 1: 	 branch_block_stmt_2486/assign_stmt_2831__exit__
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/$entry
      -- 
    cr_7335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2622_inst_req_1); -- 
    rr_7330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2622_inst_req_0); -- 
    rr_7284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2608_inst_req_0); -- 
    rr_7307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2615_inst_req_0); -- 
    rr_7353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2628_inst_req_0); -- 
    cr_7358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2628_inst_req_1); -- 
    cr_7289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2608_inst_req_1); -- 
    cr_7312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(1), ack => type_cast_2615_inst_req_1); -- 
    convTransposeD_CP_6563_elements(1) <= convTransposeD_CP_6563_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_update_start_
      -- 
    ra_6612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2488_inst_ack_0, ack => convTransposeD_CP_6563_elements(2)); -- 
    cr_6616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(2), ack => RPIPE_Block3_start_2488_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2488_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Sample/$entry
      -- 
    ca_6617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2488_inst_ack_1, ack => convTransposeD_CP_6563_elements(3)); -- 
    rr_6625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(3), ack => RPIPE_Block3_start_2491_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_update_start_
      -- 
    ra_6626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2491_inst_ack_0, ack => convTransposeD_CP_6563_elements(4)); -- 
    cr_6630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(4), ack => RPIPE_Block3_start_2491_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2491_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Sample/rr
      -- 
    ca_6631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2491_inst_ack_1, ack => convTransposeD_CP_6563_elements(5)); -- 
    rr_6639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(5), ack => RPIPE_Block3_start_2494_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Update/cr
      -- 
    ra_6640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2494_inst_ack_0, ack => convTransposeD_CP_6563_elements(6)); -- 
    cr_6644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(6), ack => RPIPE_Block3_start_2494_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2494_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Sample/rr
      -- 
    ca_6645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2494_inst_ack_1, ack => convTransposeD_CP_6563_elements(7)); -- 
    rr_6653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(7), ack => RPIPE_Block3_start_2497_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Sample/$exit
      -- 
    ra_6654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2497_inst_ack_0, ack => convTransposeD_CP_6563_elements(8)); -- 
    cr_6658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(8), ack => RPIPE_Block3_start_2497_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2497_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Sample/rr
      -- 
    ca_6659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2497_inst_ack_1, ack => convTransposeD_CP_6563_elements(9)); -- 
    rr_6667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(9), ack => RPIPE_Block3_start_2500_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Update/$entry
      -- 
    ra_6668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2500_inst_ack_0, ack => convTransposeD_CP_6563_elements(10)); -- 
    cr_6672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(10), ack => RPIPE_Block3_start_2500_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2500_Update/$exit
      -- 
    ca_6673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2500_inst_ack_1, ack => convTransposeD_CP_6563_elements(11)); -- 
    rr_6681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(11), ack => RPIPE_Block3_start_2503_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_update_start_
      -- 
    ra_6682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2503_inst_ack_0, ack => convTransposeD_CP_6563_elements(12)); -- 
    cr_6686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(12), ack => RPIPE_Block3_start_2503_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2503_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Sample/rr
      -- 
    ca_6687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2503_inst_ack_1, ack => convTransposeD_CP_6563_elements(13)); -- 
    rr_6695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(13), ack => RPIPE_Block3_start_2506_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Update/cr
      -- 
    ra_6696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2506_inst_ack_0, ack => convTransposeD_CP_6563_elements(14)); -- 
    cr_6700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(14), ack => RPIPE_Block3_start_2506_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2506_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Sample/rr
      -- 
    ca_6701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2506_inst_ack_1, ack => convTransposeD_CP_6563_elements(15)); -- 
    rr_6709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(15), ack => RPIPE_Block3_start_2509_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Update/cr
      -- 
    ra_6710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2509_inst_ack_0, ack => convTransposeD_CP_6563_elements(16)); -- 
    cr_6714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(16), ack => RPIPE_Block3_start_2509_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2509_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Sample/rr
      -- 
    ca_6715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2509_inst_ack_1, ack => convTransposeD_CP_6563_elements(17)); -- 
    rr_6723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(17), ack => RPIPE_Block3_start_2512_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Update/cr
      -- 
    ra_6724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2512_inst_ack_0, ack => convTransposeD_CP_6563_elements(18)); -- 
    cr_6728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(18), ack => RPIPE_Block3_start_2512_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2512_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Sample/rr
      -- 
    ca_6729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2512_inst_ack_1, ack => convTransposeD_CP_6563_elements(19)); -- 
    rr_6737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(19), ack => RPIPE_Block3_start_2515_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Update/cr
      -- 
    ra_6738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2515_inst_ack_0, ack => convTransposeD_CP_6563_elements(20)); -- 
    cr_6742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(20), ack => RPIPE_Block3_start_2515_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2515_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Sample/rr
      -- 
    ca_6743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2515_inst_ack_1, ack => convTransposeD_CP_6563_elements(21)); -- 
    rr_6751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(21), ack => type_cast_2519_inst_req_0); -- 
    rr_6765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(21), ack => RPIPE_Block3_start_2528_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Sample/ra
      -- 
    ra_6752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2519_inst_ack_0, ack => convTransposeD_CP_6563_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2519_Update/ca
      -- 
    ca_6757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2519_inst_ack_1, ack => convTransposeD_CP_6563_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Update/cr
      -- 
    ra_6766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2528_inst_ack_0, ack => convTransposeD_CP_6563_elements(24)); -- 
    cr_6770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(24), ack => RPIPE_Block3_start_2528_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2528_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Sample/rr
      -- 
    ca_6771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2528_inst_ack_1, ack => convTransposeD_CP_6563_elements(25)); -- 
    rr_6779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(25), ack => type_cast_2532_inst_req_0); -- 
    rr_6793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(25), ack => RPIPE_Block3_start_2540_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Sample/ra
      -- 
    ra_6780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2532_inst_ack_0, ack => convTransposeD_CP_6563_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/type_cast_2532_Update/ca
      -- 
    ca_6785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2532_inst_ack_1, ack => convTransposeD_CP_6563_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Update/cr
      -- 
    ra_6794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2540_inst_ack_0, ack => convTransposeD_CP_6563_elements(28)); -- 
    cr_6798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(28), ack => RPIPE_Block3_start_2540_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2540_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Sample/rr
      -- 
    ca_6799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2540_inst_ack_1, ack => convTransposeD_CP_6563_elements(29)); -- 
    rr_6807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(29), ack => RPIPE_Block3_start_2543_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Update/cr
      -- 
    ra_6808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2543_inst_ack_0, ack => convTransposeD_CP_6563_elements(30)); -- 
    cr_6812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(30), ack => RPIPE_Block3_start_2543_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2543_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Sample/rr
      -- 
    ca_6813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2543_inst_ack_1, ack => convTransposeD_CP_6563_elements(31)); -- 
    rr_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(31), ack => RPIPE_Block3_start_2546_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Update/cr
      -- 
    ra_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2546_inst_ack_0, ack => convTransposeD_CP_6563_elements(32)); -- 
    cr_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(32), ack => RPIPE_Block3_start_2546_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/RPIPE_Block3_start_2546_Update/ca
      -- 
    ca_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2546_inst_ack_1, ack => convTransposeD_CP_6563_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547__exit__
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599__entry__
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2489_to_assign_stmt_2547/$exit
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Update/cr
      -- 
    rr_6838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(34), ack => type_cast_2590_inst_req_0); -- 
    cr_6843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(34), ack => type_cast_2590_inst_req_1); -- 
    rr_6852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(34), ack => type_cast_2594_inst_req_0); -- 
    cr_6857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(34), ack => type_cast_2594_inst_req_1); -- 
    rr_6866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(34), ack => type_cast_2598_inst_req_0); -- 
    cr_6871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(34), ack => type_cast_2598_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(23) & convTransposeD_CP_6563_elements(27) & convTransposeD_CP_6563_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Sample/ra
      -- 
    ra_6839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2590_inst_ack_0, ack => convTransposeD_CP_6563_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2590_Update/ca
      -- 
    ca_6844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2590_inst_ack_1, ack => convTransposeD_CP_6563_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Sample/ra
      -- 
    ra_6853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2594_inst_ack_0, ack => convTransposeD_CP_6563_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2594_Update/ca
      -- 
    ca_6858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2594_inst_ack_1, ack => convTransposeD_CP_6563_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Sample/ra
      -- 
    ra_6867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_0, ack => convTransposeD_CP_6563_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/type_cast_2598_Update/ca
      -- 
    ca_6872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_1, ack => convTransposeD_CP_6563_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599__exit__
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2616/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/assign_stmt_2554_to_assign_stmt_2599/$exit
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2602/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2609/$entry
      -- CP-element group 41: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/$entry
      -- 
    rr_7258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(41), ack => type_cast_2626_inst_req_0); -- 
    cr_7263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(41), ack => type_cast_2626_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(36) & convTransposeD_CP_6563_elements(38) & convTransposeD_CP_6563_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Sample/ra
      -- 
    ra_6884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2663_inst_ack_0, ack => convTransposeD_CP_6563_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Update/ca
      -- 
    ca_6889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2663_inst_ack_1, ack => convTransposeD_CP_6563_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Sample/ra
      -- 
    ra_6898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2667_inst_ack_0, ack => convTransposeD_CP_6563_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Update/ca
      -- 
    ca_6903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2667_inst_ack_1, ack => convTransposeD_CP_6563_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Sample/ra
      -- 
    ra_6912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2671_inst_ack_0, ack => convTransposeD_CP_6563_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Update/ca
      -- 
    ca_6917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2671_inst_ack_1, ack => convTransposeD_CP_6563_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Sample/ra
      -- 
    ra_6926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2701_inst_ack_0, ack => convTransposeD_CP_6563_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Sample/req
      -- 
    ca_6931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2701_inst_ack_1, ack => convTransposeD_CP_6563_elements(49)); -- 
    req_6956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(49), ack => array_obj_ref_2707_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Sample/ack
      -- 
    ack_6957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2707_index_offset_ack_0, ack => convTransposeD_CP_6563_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_request/req
      -- 
    ack_6962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2707_index_offset_ack_1, ack => convTransposeD_CP_6563_elements(51)); -- 
    req_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(51), ack => addr_of_2708_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_request/ack
      -- 
    ack_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2708_final_reg_ack_0, ack => convTransposeD_CP_6563_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/word_access_start/word_0/rr
      -- 
    ack_6977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2708_final_reg_ack_1, ack => convTransposeD_CP_6563_elements(53)); -- 
    rr_7010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(53), ack => ptr_deref_2712_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Sample/word_access_start/word_0/ra
      -- 
    ra_7011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2712_load_0_ack_0, ack => convTransposeD_CP_6563_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/ptr_deref_2712_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/ptr_deref_2712_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/ptr_deref_2712_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/ptr_deref_2712_Merge/merge_ack
      -- 
    ca_7022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2712_load_0_ack_1, ack => convTransposeD_CP_6563_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_index_resize_1/index_resize_ack
      -- 
    req_7052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(56), ack => array_obj_ref_2730_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(43) & convTransposeD_CP_6563_elements(45) & convTransposeD_CP_6563_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_sample_complete
      -- 
    ack_7053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2730_index_offset_ack_0, ack => convTransposeD_CP_6563_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_request/req
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_offset_calculated
      -- 
    ack_7058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2730_index_offset_ack_1, ack => convTransposeD_CP_6563_elements(58)); -- 
    req_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(58), ack => addr_of_2731_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_request/ack
      -- CP-element group 59: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_sample_completed_
      -- 
    ack_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2731_final_reg_ack_0, ack => convTransposeD_CP_6563_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_word_addrgen/root_register_ack
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_update_completed_
      -- 
    ack_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2731_final_reg_ack_1, ack => convTransposeD_CP_6563_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/word_access_start/word_0/rr
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/ptr_deref_2734_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/ptr_deref_2734_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/ptr_deref_2734_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/ptr_deref_2734_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/$entry
      -- 
    rr_7111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(61), ack => ptr_deref_2734_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(55) & convTransposeD_CP_6563_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/word_access_start/word_0/ra
      -- CP-element group 62: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Sample/$exit
      -- 
    ra_7112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2734_store_0_ack_0, ack => convTransposeD_CP_6563_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/word_access_complete/word_0/ca
      -- 
    ca_7123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2734_store_0_ack_1, ack => convTransposeD_CP_6563_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Sample/ra
      -- 
    ra_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_0, ack => convTransposeD_CP_6563_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Update/$exit
      -- 
    ca_7137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_1, ack => convTransposeD_CP_6563_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751__exit__
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752__entry__
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/$exit
      -- CP-element group 66: 	 branch_block_stmt_2486/if_stmt_2752_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2486/R_cmp_2753_place
      -- 
    branch_req_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(66), ack => if_stmt_2752_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(50) & convTransposeD_CP_6563_elements(57) & convTransposeD_CP_6563_elements(63) & convTransposeD_CP_6563_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2486/merge_stmt_2758_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2486/merge_stmt_2758__exit__
      -- CP-element group 67: 	 branch_block_stmt_2486/assign_stmt_2764__entry__
      -- CP-element group 67: 	 branch_block_stmt_2486/assign_stmt_2764__exit__
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2486/if_stmt_2752_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2486/if_stmt_2752_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2486/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2486/assign_stmt_2764/$exit
      -- CP-element group 67: 	 branch_block_stmt_2486/assign_stmt_2764/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2486/merge_stmt_2758_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/merge_stmt_2758_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2486/merge_stmt_2758_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2752_branch_ack_1, ack => convTransposeD_CP_6563_elements(67)); -- 
    rr_7468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(67), ack => type_cast_2809_inst_req_0); -- 
    cr_7473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(67), ack => type_cast_2809_inst_req_1); -- 
    rr_7491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(67), ack => type_cast_2816_inst_req_0); -- 
    cr_7496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(67), ack => type_cast_2816_inst_req_1); -- 
    rr_7514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(67), ack => type_cast_2822_inst_req_0); -- 
    cr_7519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(67), ack => type_cast_2822_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2486/merge_stmt_2766_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2486/if_stmt_2752_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2486/merge_stmt_2766__exit__
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798__entry__
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2486/if_stmt_2752_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2486/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/$entry
      -- CP-element group 68: 	 branch_block_stmt_2486/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2486/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2486/merge_stmt_2766_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2486/merge_stmt_2766_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2486/merge_stmt_2766_PhiAck/dummy
      -- 
    else_choice_transition_7154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2752_branch_ack_0, ack => convTransposeD_CP_6563_elements(68)); -- 
    cr_7175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(68), ack => type_cast_2780_inst_req_1); -- 
    rr_7170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(68), ack => type_cast_2780_inst_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_sample_completed_
      -- 
    ra_7171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_0, ack => convTransposeD_CP_6563_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799_else_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798__exit__
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799__entry__
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/type_cast_2780_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2486/R_cmp121_2800_place
      -- CP-element group 70: 	 branch_block_stmt_2486/if_stmt_2799_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2486/assign_stmt_2772_to_assign_stmt_2798/$exit
      -- 
    ca_7176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_1, ack => convTransposeD_CP_6563_elements(70)); -- 
    branch_req_7184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(70), ack => if_stmt_2799_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2486/assign_stmt_2838/$entry
      -- CP-element group 71: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2486/merge_stmt_2833_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2486/if_stmt_2799_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2486/merge_stmt_2833__exit__
      -- CP-element group 71: 	 branch_block_stmt_2486/assign_stmt_2838__entry__
      -- CP-element group 71: 	 branch_block_stmt_2486/if_stmt_2799_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2486/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2486/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2486/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2486/merge_stmt_2833_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2486/merge_stmt_2833_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2486/merge_stmt_2833_PhiAck/dummy
      -- 
    if_choice_transition_7189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2799_branch_ack_1, ack => convTransposeD_CP_6563_elements(71)); -- 
    req_7209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(71), ack => WPIPE_Block3_done_2835_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2486/if_stmt_2799_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2486/if_stmt_2799_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2806/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2799_branch_ack_0, ack => convTransposeD_CP_6563_elements(72)); -- 
    rr_7419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(72), ack => type_cast_2818_inst_req_0); -- 
    cr_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(72), ack => type_cast_2818_inst_req_1); -- 
    rr_7442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(72), ack => type_cast_2824_inst_req_0); -- 
    cr_7447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(72), ack => type_cast_2824_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Update/req
      -- CP-element group 73: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_update_start_
      -- 
    ack_7210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2835_inst_ack_0, ack => convTransposeD_CP_6563_elements(73)); -- 
    req_7214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(73), ack => WPIPE_Block3_done_2835_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 branch_block_stmt_2486/assign_stmt_2838/$exit
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2486/$exit
      -- CP-element group 74: 	 branch_block_stmt_2486/branch_block_stmt_2486__exit__
      -- CP-element group 74: 	 branch_block_stmt_2486/assign_stmt_2838__exit__
      -- CP-element group 74: 	 branch_block_stmt_2486/return__
      -- CP-element group 74: 	 branch_block_stmt_2486/merge_stmt_2840__exit__
      -- CP-element group 74: 	 branch_block_stmt_2486/merge_stmt_2840_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2486/assign_stmt_2838/WPIPE_Block3_done_2835_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2486/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2486/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2486/merge_stmt_2840_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2486/merge_stmt_2840_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2486/merge_stmt_2840_PhiAck/dummy
      -- 
    ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2835_inst_ack_1, ack => convTransposeD_CP_6563_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2606_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2602/$exit
      -- CP-element group 75: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_req
      -- 
    phi_stmt_2602_req_7226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2602_req_7226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(75), ack => phi_stmt_2602_req_0); -- 
    -- Element group convTransposeD_CP_6563_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6563_elements(41), ack => convTransposeD_CP_6563_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_req
      -- CP-element group 76: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2613_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2609/$exit
      -- 
    phi_stmt_2609_req_7234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2609_req_7234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(76), ack => phi_stmt_2609_req_0); -- 
    -- Element group convTransposeD_CP_6563_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6563_elements(41), ack => convTransposeD_CP_6563_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2620_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_req
      -- CP-element group 77: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2616/$exit
      -- 
    phi_stmt_2616_req_7242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2616_req_7242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(77), ack => phi_stmt_2616_req_0); -- 
    -- Element group convTransposeD_CP_6563_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6563_elements(41), ack => convTransposeD_CP_6563_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Sample/ra
      -- 
    ra_7259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2626_inst_ack_0, ack => convTransposeD_CP_6563_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/Update/ca
      -- 
    ca_7264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2626_inst_ack_1, ack => convTransposeD_CP_6563_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_req
      -- CP-element group 80: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/$exit
      -- CP-element group 80: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2626/$exit
      -- CP-element group 80: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/$exit
      -- 
    phi_stmt_2623_req_7265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2623_req_7265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(80), ack => phi_stmt_2623_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(78) & convTransposeD_CP_6563_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2486/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(75) & convTransposeD_CP_6563_elements(76) & convTransposeD_CP_6563_elements(77) & convTransposeD_CP_6563_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Sample/ra
      -- 
    ra_7285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2608_inst_ack_0, ack => convTransposeD_CP_6563_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/ca
      -- CP-element group 83: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/Update/$exit
      -- 
    ca_7290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2608_inst_ack_1, ack => convTransposeD_CP_6563_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/$exit
      -- CP-element group 84: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/$exit
      -- CP-element group 84: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_req
      -- CP-element group 84: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2602/phi_stmt_2602_sources/type_cast_2608/SplitProtocol/$exit
      -- 
    phi_stmt_2602_req_7291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2602_req_7291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(84), ack => phi_stmt_2602_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(82) & convTransposeD_CP_6563_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Sample/ra
      -- 
    ra_7308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2615_inst_ack_0, ack => convTransposeD_CP_6563_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/Update/$exit
      -- 
    ca_7313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2615_inst_ack_1, ack => convTransposeD_CP_6563_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_req
      -- CP-element group 87: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/$exit
      -- CP-element group 87: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2609/phi_stmt_2609_sources/type_cast_2615/$exit
      -- 
    phi_stmt_2609_req_7314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2609_req_7314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(87), ack => phi_stmt_2609_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(85) & convTransposeD_CP_6563_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Sample/ra
      -- 
    ra_7331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2622_inst_ack_0, ack => convTransposeD_CP_6563_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Update/ca
      -- CP-element group 89: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/Update/$exit
      -- 
    ca_7336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2622_inst_ack_1, ack => convTransposeD_CP_6563_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/$exit
      -- CP-element group 90: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/type_cast_2622/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_req
      -- CP-element group 90: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/phi_stmt_2616_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2616/$exit
      -- 
    phi_stmt_2616_req_7337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2616_req_7337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(90), ack => phi_stmt_2616_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(88) & convTransposeD_CP_6563_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Sample/$exit
      -- 
    ra_7354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2628_inst_ack_0, ack => convTransposeD_CP_6563_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/Update/ca
      -- 
    ca_7359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2628_inst_ack_1, ack => convTransposeD_CP_6563_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/$exit
      -- CP-element group 93: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_sources/type_cast_2628/$exit
      -- CP-element group 93: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2623/phi_stmt_2623_req
      -- 
    phi_stmt_2623_req_7360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2623_req_7360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(93), ack => phi_stmt_2623_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(91) & convTransposeD_CP_6563_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2486/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(84) & convTransposeD_CP_6563_elements(87) & convTransposeD_CP_6563_elements(90) & convTransposeD_CP_6563_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2486/merge_stmt_2601_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2486/merge_stmt_2601_PhiAck/$entry
      -- 
    convTransposeD_CP_6563_elements(95) <= OrReduce(convTransposeD_CP_6563_elements(81) & convTransposeD_CP_6563_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2486/merge_stmt_2601_PhiAck/phi_stmt_2602_ack
      -- 
    phi_stmt_2602_ack_7365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2602_ack_0, ack => convTransposeD_CP_6563_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2486/merge_stmt_2601_PhiAck/phi_stmt_2609_ack
      -- 
    phi_stmt_2609_ack_7366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2609_ack_0, ack => convTransposeD_CP_6563_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2486/merge_stmt_2601_PhiAck/phi_stmt_2616_ack
      -- 
    phi_stmt_2616_ack_7367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2616_ack_0, ack => convTransposeD_CP_6563_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2486/merge_stmt_2601_PhiAck/phi_stmt_2623_ack
      -- 
    phi_stmt_2623_ack_7368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2623_ack_0, ack => convTransposeD_CP_6563_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2734_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/merge_stmt_2601_PhiAck/$exit
      -- CP-element group 100: 	 branch_block_stmt_2486/merge_stmt_2601__exit__
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751__entry__
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2663_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2667_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2671_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2739_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2730_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/type_cast_2701_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/array_obj_ref_2707_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2708_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/ptr_deref_2712_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2486/assign_stmt_2635_to_assign_stmt_2751/addr_of_2731_update_start_
      -- 
    req_7072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => addr_of_2731_final_reg_req_1); -- 
    cr_7122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => ptr_deref_2734_store_0_req_1); -- 
    rr_6883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2663_inst_req_0); -- 
    cr_6888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2663_inst_req_1); -- 
    cr_7136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2739_inst_req_1); -- 
    rr_6897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2667_inst_req_0); -- 
    cr_6902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2667_inst_req_1); -- 
    req_7057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => array_obj_ref_2730_index_offset_req_1); -- 
    rr_6911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2671_inst_req_0); -- 
    cr_6916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2671_inst_req_1); -- 
    rr_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2739_inst_req_0); -- 
    rr_6925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2701_inst_req_0); -- 
    cr_6930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => type_cast_2701_inst_req_1); -- 
    req_6961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => array_obj_ref_2707_index_offset_req_1); -- 
    req_6976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => addr_of_2708_final_reg_req_1); -- 
    cr_7021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(100), ack => ptr_deref_2712_load_0_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(96) & convTransposeD_CP_6563_elements(97) & convTransposeD_CP_6563_elements(98) & convTransposeD_CP_6563_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2806/$exit
      -- CP-element group 101: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2812_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_req
      -- 
    phi_stmt_2806_req_7403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2806_req_7403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(101), ack => phi_stmt_2806_req_1); -- 
    -- Element group convTransposeD_CP_6563_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6563_elements(72), ack => convTransposeD_CP_6563_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Sample/ra
      -- 
    ra_7420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2818_inst_ack_0, ack => convTransposeD_CP_6563_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/Update/ca
      -- 
    ca_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2818_inst_ack_1, ack => convTransposeD_CP_6563_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/$exit
      -- CP-element group 104: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/$exit
      -- CP-element group 104: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2818/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_req
      -- 
    phi_stmt_2813_req_7426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2813_req_7426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(104), ack => phi_stmt_2813_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(102) & convTransposeD_CP_6563_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Sample/ra
      -- 
    ra_7443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2824_inst_ack_0, ack => convTransposeD_CP_6563_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/Update/ca
      -- 
    ca_7448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2824_inst_ack_1, ack => convTransposeD_CP_6563_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/$exit
      -- CP-element group 107: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/$exit
      -- CP-element group 107: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2824/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_req
      -- 
    phi_stmt_2819_req_7449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2819_req_7449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(107), ack => phi_stmt_2819_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(105) & convTransposeD_CP_6563_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2486/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(101) & convTransposeD_CP_6563_elements(104) & convTransposeD_CP_6563_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Sample/ra
      -- 
    ra_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_0, ack => convTransposeD_CP_6563_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/Update/ca
      -- 
    ca_7474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_1, ack => convTransposeD_CP_6563_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/$exit
      -- CP-element group 111: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/$exit
      -- CP-element group 111: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_sources/type_cast_2809/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2806/phi_stmt_2806_req
      -- 
    phi_stmt_2806_req_7475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2806_req_7475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(111), ack => phi_stmt_2806_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(109) & convTransposeD_CP_6563_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Sample/ra
      -- 
    ra_7492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2816_inst_ack_0, ack => convTransposeD_CP_6563_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/Update/ca
      -- 
    ca_7497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2816_inst_ack_1, ack => convTransposeD_CP_6563_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/$exit
      -- CP-element group 114: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/$exit
      -- CP-element group 114: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_sources/type_cast_2816/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2813/phi_stmt_2813_req
      -- 
    phi_stmt_2813_req_7498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2813_req_7498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(114), ack => phi_stmt_2813_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(112) & convTransposeD_CP_6563_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Sample/ra
      -- 
    ra_7515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_0, ack => convTransposeD_CP_6563_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/Update/ca
      -- 
    ca_7520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_1, ack => convTransposeD_CP_6563_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/$exit
      -- CP-element group 117: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/$exit
      -- CP-element group 117: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_sources/type_cast_2822/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2819/phi_stmt_2819_req
      -- 
    phi_stmt_2819_req_7521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2819_req_7521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6563_elements(117), ack => phi_stmt_2819_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(115) & convTransposeD_CP_6563_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2486/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(111) & convTransposeD_CP_6563_elements(114) & convTransposeD_CP_6563_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2486/merge_stmt_2805_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2486/merge_stmt_2805_PhiAck/$entry
      -- 
    convTransposeD_CP_6563_elements(119) <= OrReduce(convTransposeD_CP_6563_elements(108) & convTransposeD_CP_6563_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2486/merge_stmt_2805_PhiAck/phi_stmt_2806_ack
      -- 
    phi_stmt_2806_ack_7526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2806_ack_0, ack => convTransposeD_CP_6563_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2486/merge_stmt_2805_PhiAck/phi_stmt_2813_ack
      -- 
    phi_stmt_2813_ack_7527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2813_ack_0, ack => convTransposeD_CP_6563_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2486/merge_stmt_2805_PhiAck/phi_stmt_2819_ack
      -- 
    phi_stmt_2819_ack_7528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2819_ack_0, ack => convTransposeD_CP_6563_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2486/merge_stmt_2805_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6563_elements(120) & convTransposeD_CP_6563_elements(121) & convTransposeD_CP_6563_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6563_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2729_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2729_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2706_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2706_scaled : std_logic_vector(13 downto 0);
    signal add103_2764 : std_logic_vector(15 downto 0);
    signal add32_2565 : std_logic_vector(15 downto 0);
    signal add50_2571 : std_logic_vector(15 downto 0);
    signal add63_2582 : std_logic_vector(15 downto 0);
    signal add82_2682 : std_logic_vector(63 downto 0);
    signal add84_2692 : std_logic_vector(63 downto 0);
    signal add96_2746 : std_logic_vector(31 downto 0);
    signal add_2538 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2640 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2707_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2707_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2707_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2707_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2707_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2707_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2730_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2730_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2730_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2730_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2730_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2730_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2709 : std_logic_vector(31 downto 0);
    signal arrayidx92_2732 : std_logic_vector(31 downto 0);
    signal call11_2507 : std_logic_vector(15 downto 0);
    signal call13_2510 : std_logic_vector(15 downto 0);
    signal call14_2513 : std_logic_vector(15 downto 0);
    signal call15_2516 : std_logic_vector(15 downto 0);
    signal call16_2529 : std_logic_vector(15 downto 0);
    signal call18_2541 : std_logic_vector(15 downto 0);
    signal call1_2492 : std_logic_vector(15 downto 0);
    signal call20_2544 : std_logic_vector(15 downto 0);
    signal call22_2547 : std_logic_vector(15 downto 0);
    signal call3_2495 : std_logic_vector(15 downto 0);
    signal call5_2498 : std_logic_vector(15 downto 0);
    signal call7_2501 : std_logic_vector(15 downto 0);
    signal call9_2504 : std_logic_vector(15 downto 0);
    signal call_2489 : std_logic_vector(15 downto 0);
    signal cmp111_2777 : std_logic_vector(0 downto 0);
    signal cmp121_2798 : std_logic_vector(0 downto 0);
    signal cmp_2751 : std_logic_vector(0 downto 0);
    signal conv17_2533 : std_logic_vector(31 downto 0);
    signal conv70_2664 : std_logic_vector(63 downto 0);
    signal conv73_2591 : std_logic_vector(63 downto 0);
    signal conv75_2668 : std_logic_vector(63 downto 0);
    signal conv78_2595 : std_logic_vector(63 downto 0);
    signal conv80_2672 : std_logic_vector(63 downto 0);
    signal conv95_2740 : std_logic_vector(31 downto 0);
    signal conv99_2599 : std_logic_vector(31 downto 0);
    signal conv_2520 : std_logic_vector(31 downto 0);
    signal idxprom91_2725 : std_logic_vector(63 downto 0);
    signal idxprom_2702 : std_logic_vector(63 downto 0);
    signal inc115_2781 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2786 : std_logic_vector(15 downto 0);
    signal inc_2772 : std_logic_vector(15 downto 0);
    signal indvar_2602 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2831 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2819 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2623 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2813 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2616 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2793 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2806 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2609 : std_logic_vector(15 downto 0);
    signal mul59_2655 : std_logic_vector(15 downto 0);
    signal mul81_2677 : std_logic_vector(63 downto 0);
    signal mul83_2687 : std_logic_vector(63 downto 0);
    signal mul_2645 : std_logic_vector(15 downto 0);
    signal ptr_deref_2712_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2712_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2712_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2712_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2712_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2734_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2734_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2734_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2734_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2734_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2734_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2526 : std_logic_vector(31 downto 0);
    signal shr135_2554 : std_logic_vector(15 downto 0);
    signal shr31136_2560 : std_logic_vector(15 downto 0);
    signal shr86_2698 : std_logic_vector(31 downto 0);
    signal shr90_2719 : std_logic_vector(63 downto 0);
    signal sub53_2650 : std_logic_vector(15 downto 0);
    signal sub66_2587 : std_logic_vector(15 downto 0);
    signal sub67_2660 : std_logic_vector(15 downto 0);
    signal sub_2576 : std_logic_vector(15 downto 0);
    signal tmp1_2635 : std_logic_vector(31 downto 0);
    signal tmp88_2713 : std_logic_vector(63 downto 0);
    signal type_cast_2524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2552_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2569_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2580_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2606_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2608_wire : std_logic_vector(31 downto 0);
    signal type_cast_2613_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2615_wire : std_logic_vector(15 downto 0);
    signal type_cast_2620_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2622_wire : std_logic_vector(15 downto 0);
    signal type_cast_2626_wire : std_logic_vector(15 downto 0);
    signal type_cast_2628_wire : std_logic_vector(15 downto 0);
    signal type_cast_2633_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2696_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2717_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2723_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2744_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2762_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2770_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2790_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2809_wire : std_logic_vector(15 downto 0);
    signal type_cast_2812_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2816_wire : std_logic_vector(15 downto 0);
    signal type_cast_2818_wire : std_logic_vector(15 downto 0);
    signal type_cast_2822_wire : std_logic_vector(15 downto 0);
    signal type_cast_2824_wire : std_logic_vector(15 downto 0);
    signal type_cast_2829_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2837_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2707_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2707_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2707_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2707_resized_base_address <= "00000000000000";
    array_obj_ref_2730_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2730_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2730_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2730_resized_base_address <= "00000000000000";
    ptr_deref_2712_word_offset_0 <= "00000000000000";
    ptr_deref_2734_word_offset_0 <= "00000000000000";
    type_cast_2524_wire_constant <= "00000000000000000000000000010000";
    type_cast_2552_wire_constant <= "0000000000000010";
    type_cast_2558_wire_constant <= "0000000000000001";
    type_cast_2569_wire_constant <= "1111111111111111";
    type_cast_2580_wire_constant <= "1111111111111111";
    type_cast_2606_wire_constant <= "00000000000000000000000000000000";
    type_cast_2613_wire_constant <= "0000000000000000";
    type_cast_2620_wire_constant <= "0000000000000000";
    type_cast_2633_wire_constant <= "00000000000000000000000000000100";
    type_cast_2696_wire_constant <= "00000000000000000000000000000010";
    type_cast_2717_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2723_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2744_wire_constant <= "00000000000000000000000000000100";
    type_cast_2762_wire_constant <= "0000000000000100";
    type_cast_2770_wire_constant <= "0000000000000001";
    type_cast_2790_wire_constant <= "0000000000000000";
    type_cast_2812_wire_constant <= "0000000000000000";
    type_cast_2829_wire_constant <= "00000000000000000000000000000001";
    type_cast_2837_wire_constant <= "0000000000000001";
    phi_stmt_2602: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2606_wire_constant & type_cast_2608_wire;
      req <= phi_stmt_2602_req_0 & phi_stmt_2602_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2602",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2602_ack_0,
          idata => idata,
          odata => indvar_2602,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2602
    phi_stmt_2609: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2613_wire_constant & type_cast_2615_wire;
      req <= phi_stmt_2609_req_0 & phi_stmt_2609_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2609",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2609_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2609,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2609
    phi_stmt_2616: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2620_wire_constant & type_cast_2622_wire;
      req <= phi_stmt_2616_req_0 & phi_stmt_2616_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2616",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2616_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2616,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2616
    phi_stmt_2623: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2626_wire & type_cast_2628_wire;
      req <= phi_stmt_2623_req_0 & phi_stmt_2623_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2623",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2623_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2623,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2623
    phi_stmt_2806: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2809_wire & type_cast_2812_wire_constant;
      req <= phi_stmt_2806_req_0 & phi_stmt_2806_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2806",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2806_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2806,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2806
    phi_stmt_2813: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2816_wire & type_cast_2818_wire;
      req <= phi_stmt_2813_req_0 & phi_stmt_2813_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2813",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2813_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2813,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2813
    phi_stmt_2819: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2822_wire & type_cast_2824_wire;
      req <= phi_stmt_2819_req_0 & phi_stmt_2819_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2819",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2819_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2819,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2819
    -- flow-through select operator MUX_2792_inst
    input_dim1x_x2_2793 <= type_cast_2790_wire_constant when (cmp111_2777(0) /=  '0') else inc_2772;
    addr_of_2708_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2708_final_reg_req_0;
      addr_of_2708_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2708_final_reg_req_1;
      addr_of_2708_final_reg_ack_1<= rack(0);
      addr_of_2708_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2708_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2707_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2709,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2731_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2731_final_reg_req_0;
      addr_of_2731_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2731_final_reg_req_1;
      addr_of_2731_final_reg_ack_1<= rack(0);
      addr_of_2731_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2731_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2730_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2519_inst_req_0;
      type_cast_2519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2519_inst_req_1;
      type_cast_2519_inst_ack_1<= rack(0);
      type_cast_2519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2520,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2532_inst_req_0;
      type_cast_2532_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2532_inst_req_1;
      type_cast_2532_inst_ack_1<= rack(0);
      type_cast_2532_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2532_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2533,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2590_inst_req_0;
      type_cast_2590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2590_inst_req_1;
      type_cast_2590_inst_ack_1<= rack(0);
      type_cast_2590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2594_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2594_inst_req_0;
      type_cast_2594_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2594_inst_req_1;
      type_cast_2594_inst_ack_1<= rack(0);
      type_cast_2594_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2594_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2544,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2595,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2598_inst_req_0;
      type_cast_2598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2598_inst_req_1;
      type_cast_2598_inst_ack_1<= rack(0);
      type_cast_2598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2608_inst_req_0;
      type_cast_2608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2608_inst_req_1;
      type_cast_2608_inst_ack_1<= rack(0);
      type_cast_2608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2831,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2608_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2615_inst_req_0;
      type_cast_2615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2615_inst_req_1;
      type_cast_2615_inst_ack_1<= rack(0);
      type_cast_2615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2615_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2622_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2622_inst_req_0;
      type_cast_2622_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2622_inst_req_1;
      type_cast_2622_inst_ack_1<= rack(0);
      type_cast_2622_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2622_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2813,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2622_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2626_inst_req_0;
      type_cast_2626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2626_inst_req_1;
      type_cast_2626_inst_ack_1<= rack(0);
      type_cast_2626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2626_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2628_inst_req_0;
      type_cast_2628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2628_inst_req_1;
      type_cast_2628_inst_ack_1<= rack(0);
      type_cast_2628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2628_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2628_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2663_inst_req_0;
      type_cast_2663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2663_inst_req_1;
      type_cast_2663_inst_ack_1<= rack(0);
      type_cast_2663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2609,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2667_inst_req_0;
      type_cast_2667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2667_inst_req_1;
      type_cast_2667_inst_ack_1<= rack(0);
      type_cast_2667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2667_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2668,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2671_inst_req_0;
      type_cast_2671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2671_inst_req_1;
      type_cast_2671_inst_ack_1<= rack(0);
      type_cast_2671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2650,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2701_inst_req_0;
      type_cast_2701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2701_inst_req_1;
      type_cast_2701_inst_ack_1<= rack(0);
      type_cast_2701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2739_inst_req_0;
      type_cast_2739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2739_inst_req_1;
      type_cast_2739_inst_ack_1<= rack(0);
      type_cast_2739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2609,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2780_inst_req_0;
      type_cast_2780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2780_inst_req_1;
      type_cast_2780_inst_ack_1<= rack(0);
      type_cast_2780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2781,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2809_inst_req_0;
      type_cast_2809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2809_inst_req_1;
      type_cast_2809_inst_ack_1<= rack(0);
      type_cast_2809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2809_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2816_inst_req_0;
      type_cast_2816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2816_inst_req_1;
      type_cast_2816_inst_ack_1<= rack(0);
      type_cast_2816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2616,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2816_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2818_inst_req_0;
      type_cast_2818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2818_inst_req_1;
      type_cast_2818_inst_ack_1<= rack(0);
      type_cast_2818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2818_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2818_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2822_inst_req_0;
      type_cast_2822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2822_inst_req_1;
      type_cast_2822_inst_ack_1<= rack(0);
      type_cast_2822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2824_inst_req_0;
      type_cast_2824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2824_inst_req_1;
      type_cast_2824_inst_ack_1<= rack(0);
      type_cast_2824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2824_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2707_index_1_rename
    process(R_idxprom_2706_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2706_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2706_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2707_index_1_resize
    process(idxprom_2702) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2702;
      ov := iv(13 downto 0);
      R_idxprom_2706_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2707_root_address_inst
    process(array_obj_ref_2707_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2707_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2707_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2730_index_1_rename
    process(R_idxprom91_2729_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2729_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2729_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2730_index_1_resize
    process(idxprom91_2725) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2725;
      ov := iv(13 downto 0);
      R_idxprom91_2729_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2730_root_address_inst
    process(array_obj_ref_2730_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2730_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2730_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2712_addr_0
    process(ptr_deref_2712_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2712_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2712_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2712_base_resize
    process(arrayidx87_2709) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2709;
      ov := iv(13 downto 0);
      ptr_deref_2712_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2712_gather_scatter
    process(ptr_deref_2712_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2712_data_0;
      ov(63 downto 0) := iv;
      tmp88_2713 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2712_root_address_inst
    process(ptr_deref_2712_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2712_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2712_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_addr_0
    process(ptr_deref_2734_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2734_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2734_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_base_resize
    process(arrayidx92_2732) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2732;
      ov := iv(13 downto 0);
      ptr_deref_2734_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_gather_scatter
    process(tmp88_2713) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2713;
      ov(63 downto 0) := iv;
      ptr_deref_2734_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2734_root_address_inst
    process(ptr_deref_2734_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2734_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2734_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2752_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2751;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2752_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2752_branch_req_0,
          ack0 => if_stmt_2752_branch_ack_0,
          ack1 => if_stmt_2752_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2799_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2798;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2799_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2799_branch_req_0,
          ack0 => if_stmt_2799_branch_ack_0,
          ack1 => if_stmt_2799_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2564_inst
    process(shr135_2554, shr31136_2560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2554, shr31136_2560, tmp_var);
      add32_2565 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2570_inst
    process(call7_2501) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2501, type_cast_2569_wire_constant, tmp_var);
      add50_2571 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2581_inst
    process(call9_2504) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2504, type_cast_2580_wire_constant, tmp_var);
      add63_2582 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2649_inst
    process(sub_2576, mul_2645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2576, mul_2645, tmp_var);
      sub53_2650 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2659_inst
    process(sub66_2587, mul59_2655) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2587, mul59_2655, tmp_var);
      sub67_2660 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2763_inst
    process(input_dim2x_x1_2609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2609, type_cast_2762_wire_constant, tmp_var);
      add103_2764 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2771_inst
    process(input_dim1x_x1_2616) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2616, type_cast_2770_wire_constant, tmp_var);
      inc_2772 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2785_inst
    process(inc115_2781, input_dim0x_x2_2623) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2781, input_dim0x_x2_2623, tmp_var);
      inc115x_xinput_dim0x_x2_2786 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2639_inst
    process(add_2538, tmp1_2635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2538, tmp1_2635, tmp_var);
      add_src_0x_x0_2640 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2745_inst
    process(conv95_2740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2740, type_cast_2744_wire_constant, tmp_var);
      add96_2746 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2830_inst
    process(indvar_2602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2602, type_cast_2829_wire_constant, tmp_var);
      indvarx_xnext_2831 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2681_inst
    process(mul81_2677, conv75_2668) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2677, conv75_2668, tmp_var);
      add82_2682 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2691_inst
    process(mul83_2687, conv70_2664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2687, conv70_2664, tmp_var);
      add84_2692 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2724_inst
    process(shr90_2719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2719, type_cast_2723_wire_constant, tmp_var);
      idxprom91_2725 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2776_inst
    process(inc_2772, call1_2492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2772, call1_2492, tmp_var);
      cmp111_2777 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2797_inst
    process(inc115x_xinput_dim0x_x2_2786, call_2489) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2786, call_2489, tmp_var);
      cmp121_2798 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2553_inst
    process(call_2489) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2489, type_cast_2552_wire_constant, tmp_var);
      shr135_2554 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2559_inst
    process(call_2489) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2489, type_cast_2558_wire_constant, tmp_var);
      shr31136_2560 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2697_inst
    process(add_src_0x_x0_2640) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2640, type_cast_2696_wire_constant, tmp_var);
      shr86_2698 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2718_inst
    process(add84_2692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2692, type_cast_2717_wire_constant, tmp_var);
      shr90_2719 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2644_inst
    process(input_dim0x_x2_2623, call13_2510) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2623, call13_2510, tmp_var);
      mul_2645 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2654_inst
    process(input_dim1x_x1_2616, call13_2510) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2616, call13_2510, tmp_var);
      mul59_2655 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2634_inst
    process(indvar_2602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2602, type_cast_2633_wire_constant, tmp_var);
      tmp1_2635 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2676_inst
    process(conv80_2672, conv78_2595) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2672, conv78_2595, tmp_var);
      mul81_2677 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2686_inst
    process(add82_2682, conv73_2591) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2682, conv73_2591, tmp_var);
      mul83_2687 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2537_inst
    process(shl_2526, conv17_2533) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2526, conv17_2533, tmp_var);
      add_2538 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2525_inst
    process(conv_2520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2520, type_cast_2524_wire_constant, tmp_var);
      shl_2526 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2575_inst
    process(add50_2571, call14_2513) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2571, call14_2513, tmp_var);
      sub_2576 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2586_inst
    process(add63_2582, call14_2513) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2582, call14_2513, tmp_var);
      sub66_2587 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2750_inst
    process(add96_2746, conv99_2599) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2746, conv99_2599, tmp_var);
      cmp_2751 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2707_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2706_scaled;
      array_obj_ref_2707_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2707_index_offset_req_0;
      array_obj_ref_2707_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2707_index_offset_req_1;
      array_obj_ref_2707_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2730_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2729_scaled;
      array_obj_ref_2730_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2730_index_offset_req_0;
      array_obj_ref_2730_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2730_index_offset_req_1;
      array_obj_ref_2730_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2712_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2712_load_0_req_0;
      ptr_deref_2712_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2712_load_0_req_1;
      ptr_deref_2712_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2712_word_address_0;
      ptr_deref_2712_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2734_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2734_store_0_req_0;
      ptr_deref_2734_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2734_store_0_req_1;
      ptr_deref_2734_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2734_word_address_0;
      data_in <= ptr_deref_2734_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2488_inst RPIPE_Block3_start_2491_inst RPIPE_Block3_start_2494_inst RPIPE_Block3_start_2497_inst RPIPE_Block3_start_2500_inst RPIPE_Block3_start_2503_inst RPIPE_Block3_start_2506_inst RPIPE_Block3_start_2509_inst RPIPE_Block3_start_2512_inst RPIPE_Block3_start_2515_inst RPIPE_Block3_start_2528_inst RPIPE_Block3_start_2540_inst RPIPE_Block3_start_2543_inst RPIPE_Block3_start_2546_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2488_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2491_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2494_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2497_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2500_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2503_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2506_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2509_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2512_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2515_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2528_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2540_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2543_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2546_inst_req_0;
      RPIPE_Block3_start_2488_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2491_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2494_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2497_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2500_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2503_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2506_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2509_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2512_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2515_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2528_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2540_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2543_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2546_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2488_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2491_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2494_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2497_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2500_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2503_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2506_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2509_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2512_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2515_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2528_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2540_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2543_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2546_inst_req_1;
      RPIPE_Block3_start_2488_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2491_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2494_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2497_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2500_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2503_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2506_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2509_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2512_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2515_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2528_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2540_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2543_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2546_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2489 <= data_out(223 downto 208);
      call1_2492 <= data_out(207 downto 192);
      call3_2495 <= data_out(191 downto 176);
      call5_2498 <= data_out(175 downto 160);
      call7_2501 <= data_out(159 downto 144);
      call9_2504 <= data_out(143 downto 128);
      call11_2507 <= data_out(127 downto 112);
      call13_2510 <= data_out(111 downto 96);
      call14_2513 <= data_out(95 downto 80);
      call15_2516 <= data_out(79 downto 64);
      call16_2529 <= data_out(63 downto 48);
      call18_2541 <= data_out(47 downto 32);
      call20_2544 <= data_out(31 downto 16);
      call22_2547 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2835_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2835_inst_req_0;
      WPIPE_Block3_done_2835_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2835_inst_req_1;
      WPIPE_Block3_done_2835_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2837_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_29_load_0_req_0 : boolean;
  signal LOAD_count_29_load_0_ack_0 : boolean;
  signal LOAD_count_29_load_0_req_1 : boolean;
  signal LOAD_count_29_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_30/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_update_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/$entry
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$entry
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_30/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_29_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_29_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_29_word_address_0 <= "0";
    -- equivalence LOAD_count_29_gather_scatter
    process(LOAD_count_29_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_29_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_29_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_29_load_0_req_0;
      LOAD_count_29_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_29_load_0_req_1;
      LOAD_count_29_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_29_word_address_0;
      LOAD_count_29_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
