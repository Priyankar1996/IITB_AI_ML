-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_44_branch_req_0 : boolean;
  signal phi_stmt_46_ack_0 : boolean;
  signal phi_stmt_46_req_1 : boolean;
  signal phi_stmt_46_req_0 : boolean;
  signal n_address_280_50_buf_req_0 : boolean;
  signal n_address_280_50_buf_ack_0 : boolean;
  signal n_address_280_50_buf_req_1 : boolean;
  signal n_address_280_50_buf_ack_1 : boolean;
  signal phi_stmt_51_req_1 : boolean;
  signal phi_stmt_51_req_0 : boolean;
  signal phi_stmt_51_ack_0 : boolean;
  signal n_word_start_269_56_buf_req_0 : boolean;
  signal n_word_start_269_56_buf_ack_0 : boolean;
  signal n_word_start_269_56_buf_req_1 : boolean;
  signal n_word_start_269_56_buf_ack_1 : boolean;
  signal n_winr_209_70_buf_req_0 : boolean;
  signal n_winr_209_70_buf_ack_0 : boolean;
  signal phi_stmt_57_req_1 : boolean;
  signal phi_stmt_57_req_0 : boolean;
  signal phi_stmt_57_ack_0 : boolean;
  signal nl_start_35_59_buf_req_0 : boolean;
  signal nl_start_35_59_buf_ack_0 : boolean;
  signal nl_start_35_59_buf_req_1 : boolean;
  signal nl_start_35_59_buf_ack_1 : boolean;
  signal n_left_288_60_buf_req_0 : boolean;
  signal n_left_288_60_buf_ack_0 : boolean;
  signal n_left_288_60_buf_req_1 : boolean;
  signal n_left_288_60_buf_ack_1 : boolean;
  signal phi_stmt_61_req_1 : boolean;
  signal phi_stmt_61_req_0 : boolean;
  signal phi_stmt_61_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal n_blk_308_65_buf_req_0 : boolean;
  signal n_blk_308_65_buf_ack_0 : boolean;
  signal n_blk_308_65_buf_req_1 : boolean;
  signal n_blk_308_65_buf_ack_1 : boolean;
  signal phi_stmt_66_req_1 : boolean;
  signal phi_stmt_66_req_0 : boolean;
  signal phi_stmt_66_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_1 : boolean;
  signal n_winr_209_70_buf_req_1 : boolean;
  signal n_winr_209_70_buf_ack_1 : boolean;
  signal phi_stmt_71_req_1 : boolean;
  signal phi_stmt_71_req_0 : boolean;
  signal phi_stmt_71_ack_0 : boolean;
  signal n_col_222_75_buf_req_0 : boolean;
  signal n_col_222_75_buf_ack_0 : boolean;
  signal n_col_222_75_buf_req_1 : boolean;
  signal n_col_222_75_buf_ack_1 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal n_row_234_78_buf_req_0 : boolean;
  signal n_row_234_78_buf_ack_0 : boolean;
  signal n_row_234_78_buf_req_1 : boolean;
  signal n_row_234_78_buf_ack_1 : boolean;
  signal array_obj_ref_133_index_offset_req_0 : boolean;
  signal array_obj_ref_133_index_offset_ack_0 : boolean;
  signal array_obj_ref_133_index_offset_req_1 : boolean;
  signal array_obj_ref_133_index_offset_ack_1 : boolean;
  signal addr_of_134_final_reg_req_0 : boolean;
  signal addr_of_134_final_reg_ack_0 : boolean;
  signal addr_of_134_final_reg_req_1 : boolean;
  signal addr_of_134_final_reg_ack_1 : boolean;
  signal ptr_deref_138_load_0_req_0 : boolean;
  signal ptr_deref_138_load_0_ack_0 : boolean;
  signal ptr_deref_138_load_0_req_1 : boolean;
  signal ptr_deref_138_load_0_ack_1 : boolean;
  signal slice_142_inst_req_0 : boolean;
  signal slice_142_inst_ack_0 : boolean;
  signal slice_142_inst_req_1 : boolean;
  signal slice_142_inst_ack_1 : boolean;
  signal slice_146_inst_req_0 : boolean;
  signal slice_146_inst_ack_0 : boolean;
  signal slice_146_inst_req_1 : boolean;
  signal slice_146_inst_ack_1 : boolean;
  signal slice_150_inst_req_0 : boolean;
  signal slice_150_inst_ack_0 : boolean;
  signal slice_150_inst_req_1 : boolean;
  signal slice_150_inst_ack_1 : boolean;
  signal slice_154_inst_req_0 : boolean;
  signal slice_154_inst_ack_0 : boolean;
  signal slice_154_inst_req_1 : boolean;
  signal slice_154_inst_ack_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_1 : boolean;
  signal do_while_stmt_44_branch_ack_0 : boolean;
  signal do_while_stmt_44_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__exit__
      -- CP-element group 0: 	 branch_block_stmt_26/do_while_stmt_44__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_26/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/branch_block_stmt_26__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_26/$exit
      -- CP-element group 1: 	 branch_block_stmt_26/branch_block_stmt_26__exit__
      -- CP-element group 1: 	 branch_block_stmt_26/do_while_stmt_44__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/$entry
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_26/do_while_stmt_44/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/condition_done
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_26/do_while_stmt_44/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	97 
    -- CP-element group 7: 	116 
    -- CP-element group 7: 	135 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	99 
    -- CP-element group 8: 	118 
    -- CP-element group 8: 	137 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	91 
    -- CP-element group 9: 	92 
    -- CP-element group 9: 	110 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	130 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	203 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_44_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(14) & access_T_CP_0_elements(203);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	129 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	112 
    -- CP-element group 11: 	131 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(15) & access_T_CP_0_elements(32) & access_T_CP_0_elements(51) & access_T_CP_0_elements(70) & access_T_CP_0_elements(91) & access_T_CP_0_elements(110) & access_T_CP_0_elements(129) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	94 
    -- CP-element group 12: 	113 
    -- CP-element group 12: 	132 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12: 	91 
    -- CP-element group 12: 	110 
    -- CP-element group 12: 	129 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(17) & access_T_CP_0_elements(35) & access_T_CP_0_elements(54) & access_T_CP_0_elements(73) & access_T_CP_0_elements(94) & access_T_CP_0_elements(113) & access_T_CP_0_elements(132);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: 	92 
    -- CP-element group 13: 	111 
    -- CP-element group 13: 	130 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	95 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	133 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(16) & access_T_CP_0_elements(33) & access_T_CP_0_elements(52) & access_T_CP_0_elements(71) & access_T_CP_0_elements(92) & access_T_CP_0_elements(111) & access_T_CP_0_elements(130);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	96 
    -- CP-element group 14: 	115 
    -- CP-element group 14: 	134 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(56) & access_T_CP_0_elements(75) & access_T_CP_0_elements(96) & access_T_CP_0_elements(115) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	151 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (15) 
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(18), ack => array_obj_ref_133_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_trigger
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req_ps
      -- 
    phi_stmt_46_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => phi_stmt_46_req_1); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req_ps
      -- 
    phi_stmt_46_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_46_req_0); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack_ps
      -- 
    phi_stmt_46_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_46_ack_0, ack => access_T_CP_0_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start_
      -- 
    -- Element group access_T_CP_0_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed__ps
      -- 
    access_T_CP_0_elements(26) <= access_T_CP_0_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(25), ack => access_T_CP_0_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(28), ack => n_address_280_50_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_start_
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/req
      -- 
    req_76_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_76_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(29), ack => n_address_280_50_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_50_buf_ack_0, ack => access_T_CP_0_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/ack
      -- 
    ack_77_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_50_buf_ack_1, ack => access_T_CP_0_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start_
      -- 
    access_T_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	177 
    -- CP-element group 33: 	191 
    -- CP-element group 33: 	184 
    -- CP-element group 33: 	198 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start_
      -- 
    access_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(177) & access_T_CP_0_elements(191) & access_T_CP_0_elements(184) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start__ps
      -- 
    access_T_CP_0_elements(34) <= access_T_CP_0_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	196 
    -- CP-element group 37: 	175 
    -- CP-element group 37: 	189 
    -- CP-element group 37: 	182 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_trigger
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req_ps
      -- 
    phi_stmt_51_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(39), ack => phi_stmt_51_req_1); -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req_ps
      -- 
    phi_stmt_51_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_51_req_0); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack_ps
      -- 
    phi_stmt_51_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_51_ack_0, ack => access_T_CP_0_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_start_
      -- 
    -- Element group access_T_CP_0_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_completed__ps
      -- 
    access_T_CP_0_elements(45) <= access_T_CP_0_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(44), ack => access_T_CP_0_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(47), ack => n_word_start_269_56_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_start_
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/req
      -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(48), ack => n_word_start_269_56_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_56_buf_ack_0, ack => access_T_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_56_buf_ack_1, ack => access_T_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start_
      -- 
    access_T_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start_
      -- 
    access_T_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start__ps
      -- 
    access_T_CP_0_elements(53) <= access_T_CP_0_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_trigger
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req_ps
      -- 
    phi_stmt_57_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(58), ack => phi_stmt_57_req_1); -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_trigger
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req_ps
      -- 
    phi_stmt_57_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_57_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack_ps
      -- 
    phi_stmt_57_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_57_ack_0, ack => access_T_CP_0_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => nl_start_35_59_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start_
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(63), ack => nl_start_35_59_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_0, ack => access_T_CP_0_elements(64)); -- 
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_1, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(66), ack => n_left_288_60_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start_
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => n_left_288_60_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_0, ack => access_T_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_1, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start_
      -- 
    access_T_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	191 
    -- CP-element group 71: 	184 
    -- CP-element group 71: 	198 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start_
      -- 
    access_T_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(191) & access_T_CP_0_elements(184) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start__ps
      -- 
    access_T_CP_0_elements(72) <= access_T_CP_0_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	196 
    -- CP-element group 75: 	189 
    -- CP-element group 75: 	182 
    -- CP-element group 75: 	14 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_trigger
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req_ps
      -- 
    phi_stmt_61_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(77), ack => phi_stmt_61_req_1); -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req_ps
      -- 
    phi_stmt_61_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_61_req_0); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack_ps
      -- 
    phi_stmt_61_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_61_ack_0, ack => access_T_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/rr
      -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => type_cast_64_inst_req_0); -- 
    access_T_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(85);
      gj_access_T_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start_
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/cr
      -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => type_cast_64_inst_req_1); -- 
    access_T_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(82) & access_T_CP_0_elements(86);
      gj_access_T_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => access_T_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/req
      -- 
    req_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => n_blk_308_65_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start_
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/req
      -- 
    req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => n_blk_308_65_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/ack
      -- 
    ack_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/ack
      -- 
    ack_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	9 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	12 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	11 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start_
      -- 
    access_T_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	9 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	96 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	13 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start_
      -- 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(96);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	11 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start__ps
      -- 
    access_T_CP_0_elements(93) <= access_T_CP_0_elements(11);
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	12 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	13 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(13);
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	14 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	7 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_trigger
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(7);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req_ps
      -- 
    phi_stmt_66_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_66_req_1); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	8 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(8);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req_ps
      -- 
    phi_stmt_66_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_66_req_0); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack_ps
      -- 
    phi_stmt_66_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_66_ack_0, ack => access_T_CP_0_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_sample_start__ps
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_update_start__ps
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_update_start_
      -- 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_update_completed__ps
      -- 
    access_T_CP_0_elements(104) <= access_T_CP_0_elements(105);
    -- CP-element group 105:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	104 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_69_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(103), ack => access_T_CP_0_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Sample/req
      -- 
    req_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(106), ack => n_winr_209_70_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_update_start_
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Update/req
      -- 
    req_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(107), ack => n_winr_209_70_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Sample/ack
      -- 
    ack_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_70_buf_ack_0, ack => access_T_CP_0_elements(108)); -- 
    -- CP-element group 109:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_update_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_70_Update/ack
      -- 
    ack_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_70_buf_ack_1, ack => access_T_CP_0_elements(109)); -- 
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	9 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	12 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	11 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start_
      -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	115 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	13 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start_
      -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	11 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start__ps
      -- 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(11);
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	12 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(13);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	111 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	7 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(7);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req_ps
      -- 
    phi_stmt_71_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_71_req_1); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	8 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(8);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req_ps
      -- 
    phi_stmt_71_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_71_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack_ps
      -- 
    phi_stmt_71_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_71_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_start_
      -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_completed__ps
      -- 
    access_T_CP_0_elements(123) <= access_T_CP_0_elements(124);
    -- CP-element group 124:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_74_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(124) is a control-delay.
    cp_element_124_delay: control_delay_element  generic map(name => " 124_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(122), ack => access_T_CP_0_elements(124), clk => clk, reset =>reset);
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/req
      -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => n_col_222_75_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_start_
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/req
      -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(126), ack => n_col_222_75_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Sample/ack
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_75_buf_ack_0, ack => access_T_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_75_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_75_buf_ack_1, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	12 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	11 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start_
      -- 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	134 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	13 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	11 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(11);
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start__ps
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	130 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_76_req_0); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_76_req_1); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/req
      -- 
    req_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(140), ack => n_row_234_78_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_start_
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/req
      -- 
    req_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(141), ack => n_row_234_78_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Sample/ack
      -- 
    ack_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_78_buf_ack_0, ack => access_T_CP_0_elements(142)); -- 
    -- CP-element group 143:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_completed__ps
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_78_Update/ack
      -- 
    ack_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_78_buf_ack_1, ack => access_T_CP_0_elements(143)); -- 
    -- CP-element group 144:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_start_
      -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_completed__ps
      -- 
    access_T_CP_0_elements(146) <= access_T_CP_0_elements(147);
    -- CP-element group 147:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_80_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(147) is a control-delay.
    cp_element_147_delay: control_delay_element  generic map(name => " 147_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(145), ack => access_T_CP_0_elements(147), clk => clk, reset =>reset);
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_134_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_start_
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_134_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_133_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	18 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_138_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	173 
    -- CP-element group 156: 	169 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_start_
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_138_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(161) & access_T_CP_0_elements(165) & access_T_CP_0_elements(173) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	167 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	171 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_142_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_start_
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_142_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_146_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_start_
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_146_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	156 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_150_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_start_
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_150_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	156 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_154_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_start_
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_154_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	156 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	37 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_156_delayed_14_0_156_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_start_
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_156_delayed_14_0_156_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	33 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	162 
    -- CP-element group 179: 	178 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_160_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(162) & access_T_CP_0_elements(178) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: 	160 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_start_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_160_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	37 
    -- CP-element group 182: 	75 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_160_delayed_14_0_163_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_start_
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_160_delayed_14_0_163_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	33 
    -- CP-element group 184: 	71 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	166 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_167_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(185) & access_T_CP_0_elements(181) & access_T_CP_0_elements(166) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	164 
    -- CP-element group 187: 	183 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/req
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_start_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$exit
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_167_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	37 
    -- CP-element group 189: 	75 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_164_delayed_14_0_170_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_start_
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_164_delayed_14_0_170_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	33 
    -- CP-element group 191: 	71 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	170 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_174_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(188) & access_T_CP_0_elements(192) & access_T_CP_0_elements(170) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	168 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_start_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_174_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	37 
    -- CP-element group 196: 	75 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_168_delayed_14_0_177_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(37) & access_T_CP_0_elements(75) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_start_
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_168_delayed_14_0_177_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	33 
    -- CP-element group 198: 	71 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	174 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_181_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(195) & access_T_CP_0_elements(174) & access_T_CP_0_elements(199) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	172 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_start_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_181_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	179 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	151 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(151) & access_T_CP_0_elements(12) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_26/do_while_stmt_44/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_44_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_44_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_46_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(24);
      access_T_CP_0_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(19);
      access_T_CP_0_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(30);
      access_T_CP_0_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(31);
      access_T_CP_0_elements(20) <= phi_mux_reqs(1);
      phi_stmt_46_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_46_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(17), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(18), 
          phi_mux_ack => access_T_CP_0_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_51_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(43);
      access_T_CP_0_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(38);
      access_T_CP_0_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(49);
      access_T_CP_0_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(50);
      access_T_CP_0_elements(39) <= phi_mux_reqs(1);
      phi_stmt_51_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_51_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(34), 
          phi_sample_ack => access_T_CP_0_elements(35), 
          phi_update_req => access_T_CP_0_elements(36), 
          phi_update_ack => access_T_CP_0_elements(37), 
          phi_mux_ack => access_T_CP_0_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_57_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(64);
      access_T_CP_0_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(65);
      access_T_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(57);
      access_T_CP_0_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(58) <= phi_mux_reqs(1);
      phi_stmt_57_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_57_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(53), 
          phi_sample_ack => access_T_CP_0_elements(54), 
          phi_update_req => access_T_CP_0_elements(55), 
          phi_update_ack => access_T_CP_0_elements(56), 
          phi_mux_ack => access_T_CP_0_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_61_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(85);
      access_T_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(76);
      access_T_CP_0_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(77) <= phi_mux_reqs(1);
      phi_stmt_61_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_61_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(72), 
          phi_sample_ack => access_T_CP_0_elements(73), 
          phi_update_req => access_T_CP_0_elements(74), 
          phi_update_ack => access_T_CP_0_elements(75), 
          phi_mux_ack => access_T_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_66_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(102);
      access_T_CP_0_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(100) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(106)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(108);
      access_T_CP_0_elements(107)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(109);
      access_T_CP_0_elements(98) <= phi_mux_reqs(1);
      phi_stmt_66_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_66_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(93), 
          phi_sample_ack => access_T_CP_0_elements(94), 
          phi_update_req => access_T_CP_0_elements(95), 
          phi_update_ack => access_T_CP_0_elements(96), 
          phi_mux_ack => access_T_CP_0_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_71_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(121);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(119) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(117) <= phi_mux_reqs(1);
      phi_stmt_71_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_71_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(112), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(136) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(138) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_76_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(131), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_125_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_205_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_218_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_231_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_293_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_278_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_107_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_114_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_213_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_227_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_94_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_260_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_103_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_110_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_117_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_90_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_97_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_274_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_240_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_30_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_249_wire : std_logic_vector(31 downto 0);
    signal MUX_206_wire : std_logic_vector(15 downto 0);
    signal MUX_219_wire : std_logic_vector(15 downto 0);
    signal MUX_300_wire : std_logic_vector(15 downto 0);
    signal MUX_306_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_312_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_118_wire : std_logic_vector(0 downto 0);
    signal R_address_132_resized : std_logic_vector(13 downto 0);
    signal R_address_132_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_286_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_298_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_106_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_113_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_295_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_93_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_303_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_39_wire : std_logic_vector(0 downto 0);
    signal address_46 : std_logic_vector(63 downto 0);
    signal array_obj_ref_133_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_root_address : std_logic_vector(13 downto 0);
    signal c1_156_delayed_14_0_158 : std_logic_vector(0 downto 0);
    signal c1_86 : std_logic_vector(0 downto 0);
    signal c2_160_delayed_14_0_165 : std_logic_vector(0 downto 0);
    signal c2_99 : std_logic_vector(0 downto 0);
    signal c3_120 : std_logic_vector(0 downto 0);
    signal c3_164_delayed_14_0_172 : std_logic_vector(0 downto 0);
    signal c4_128 : std_logic_vector(0 downto 0);
    signal c4_168_delayed_14_0_179 : std_logic_vector(0 downto 0);
    signal col_71 : std_logic_vector(15 downto 0);
    signal col_done_198 : std_logic_vector(0 downto 0);
    signal fetch_addr_135 : std_logic_vector(31 downto 0);
    signal flag1_188 : std_logic_vector(0 downto 0);
    signal fn_blk_43 : std_logic_vector(15 downto 0);
    signal konst_102_wire_constant : std_logic_vector(1 downto 0);
    signal konst_105_wire_constant : std_logic_vector(15 downto 0);
    signal konst_109_wire_constant : std_logic_vector(1 downto 0);
    signal konst_112_wire_constant : std_logic_vector(15 downto 0);
    signal konst_116_wire_constant : std_logic_vector(1 downto 0);
    signal konst_126_wire_constant : std_logic_vector(15 downto 0);
    signal konst_202_wire_constant : std_logic_vector(15 downto 0);
    signal konst_204_wire_constant : std_logic_vector(15 downto 0);
    signal konst_215_wire_constant : std_logic_vector(15 downto 0);
    signal konst_217_wire_constant : std_logic_vector(15 downto 0);
    signal konst_230_wire_constant : std_logic_vector(15 downto 0);
    signal konst_259_wire_constant : std_logic_vector(31 downto 0);
    signal konst_267_wire_constant : std_logic_vector(1 downto 0);
    signal konst_273_wire_constant : std_logic_vector(31 downto 0);
    signal konst_277_wire_constant : std_logic_vector(63 downto 0);
    signal konst_294_wire_constant : std_logic_vector(15 downto 0);
    signal konst_296_wire_constant : std_logic_vector(15 downto 0);
    signal konst_302_wire_constant : std_logic_vector(15 downto 0);
    signal konst_305_wire_constant : std_logic_vector(15 downto 0);
    signal konst_38_wire_constant : std_logic_vector(15 downto 0);
    signal konst_41_wire_constant : std_logic_vector(15 downto 0);
    signal konst_84_wire_constant : std_logic_vector(1 downto 0);
    signal konst_89_wire_constant : std_logic_vector(1 downto 0);
    signal konst_92_wire_constant : std_logic_vector(15 downto 0);
    signal konst_96_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_32 : std_logic_vector(31 downto 0);
    signal n_address_280 : std_logic_vector(63 downto 0);
    signal n_address_280_50_buffered : std_logic_vector(63 downto 0);
    signal n_blk_308 : std_logic_vector(15 downto 0);
    signal n_blk_308_65_buffered : std_logic_vector(15 downto 0);
    signal n_col_222 : std_logic_vector(15 downto 0);
    signal n_col_222_75_buffered : std_logic_vector(15 downto 0);
    signal n_left_288 : std_logic_vector(15 downto 0);
    signal n_left_288_60_buffered : std_logic_vector(15 downto 0);
    signal n_row_234 : std_logic_vector(15 downto 0);
    signal n_row_234_78_buffered : std_logic_vector(15 downto 0);
    signal n_winr_209 : std_logic_vector(15 downto 0);
    signal n_winr_209_70_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_269 : std_logic_vector(1 downto 0);
    signal n_word_start_269_56_buffered : std_logic_vector(1 downto 0);
    signal na1_244 : std_logic_vector(31 downto 0);
    signal na2_251 : std_logic_vector(31 downto 0);
    signal na3_256 : std_logic_vector(31 downto 0);
    signal na4_262 : std_logic_vector(15 downto 0);
    signal nl_start_35 : std_logic_vector(15 downto 0);
    signal nl_start_35_59_buffered : std_logic_vector(15 downto 0);
    signal num_blk_61 : std_logic_vector(15 downto 0);
    signal num_left_57 : std_logic_vector(15 downto 0);
    signal ptr_deref_138_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_138_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_76 : std_logic_vector(15 downto 0);
    signal type_cast_124_wire : std_logic_vector(15 downto 0);
    signal type_cast_248_wire : std_logic_vector(31 downto 0);
    signal type_cast_266_wire : std_logic_vector(1 downto 0);
    signal type_cast_275_wire : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_64_wire : std_logic_vector(15 downto 0);
    signal type_cast_69_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_74_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_80_wire_constant : std_logic_vector(15 downto 0);
    signal w1_143 : std_logic_vector(15 downto 0);
    signal w2_147 : std_logic_vector(15 downto 0);
    signal w3_151 : std_logic_vector(15 downto 0);
    signal w4_155 : std_logic_vector(15 downto 0);
    signal winr_66 : std_logic_vector(15 downto 0);
    signal winr_done_193 : std_logic_vector(0 downto 0);
    signal word_read_139 : std_logic_vector(63 downto 0);
    signal word_start_51 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_133_constant_part_of_offset <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_133_resized_base_address <= "00000000000000";
    konst_102_wire_constant <= "00";
    konst_105_wire_constant <= "0000000000000010";
    konst_109_wire_constant <= "01";
    konst_112_wire_constant <= "0000000000000001";
    konst_116_wire_constant <= "10";
    konst_126_wire_constant <= "0000000000000011";
    konst_202_wire_constant <= "0000000000000000";
    konst_204_wire_constant <= "0000000000000001";
    konst_215_wire_constant <= "0000000000000000";
    konst_217_wire_constant <= "0000000000000001";
    konst_230_wire_constant <= "0000000000000001";
    konst_259_wire_constant <= "00000000000000000000000000000011";
    konst_267_wire_constant <= "00";
    konst_273_wire_constant <= "00000000000000000000000000000010";
    konst_277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_294_wire_constant <= "0000000000000100";
    konst_296_wire_constant <= "0000000000000100";
    konst_302_wire_constant <= "0000000000000100";
    konst_305_wire_constant <= "0000000000000100";
    konst_38_wire_constant <= "0000000000000100";
    konst_41_wire_constant <= "0000000000000100";
    konst_84_wire_constant <= "00";
    konst_89_wire_constant <= "00";
    konst_92_wire_constant <= "0000000000000001";
    konst_96_wire_constant <= "01";
    ptr_deref_138_word_offset_0 <= "00000000000000";
    type_cast_49_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_55_wire_constant <= "00";
    type_cast_69_wire_constant <= "0000000000000000";
    type_cast_74_wire_constant <= "0000000000000000";
    type_cast_80_wire_constant <= "0000000000000000";
    phi_stmt_46: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_49_wire_constant & n_address_280_50_buffered;
      req <= phi_stmt_46_req_0 & phi_stmt_46_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_46",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_46_ack_0,
          idata => idata,
          odata => address_46,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_46
    phi_stmt_51: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_55_wire_constant & n_word_start_269_56_buffered;
      req <= phi_stmt_51_req_0 & phi_stmt_51_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_51",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_51_ack_0,
          idata => idata,
          odata => word_start_51,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_51
    phi_stmt_57: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nl_start_35_59_buffered & n_left_288_60_buffered;
      req <= phi_stmt_57_req_0 & phi_stmt_57_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_57",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_57_ack_0,
          idata => idata,
          odata => num_left_57,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_57
    phi_stmt_61: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_64_wire & n_blk_308_65_buffered;
      req <= phi_stmt_61_req_0 & phi_stmt_61_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_61",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_61_ack_0,
          idata => idata,
          odata => num_blk_61,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_61
    phi_stmt_66: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_69_wire_constant & n_winr_209_70_buffered;
      req <= phi_stmt_66_req_0 & phi_stmt_66_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_66",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_66_ack_0,
          idata => idata,
          odata => winr_66,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_66
    phi_stmt_71: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_74_wire_constant & n_col_222_75_buffered;
      req <= phi_stmt_71_req_0 & phi_stmt_71_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_71",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_71_ack_0,
          idata => idata,
          odata => col_71,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_71
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row_234_78_buffered & type_cast_80_wire_constant;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => row_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    -- flow-through select operator MUX_206_inst
    MUX_206_wire <= konst_202_wire_constant when (winr_done_193(0) /=  '0') else ADD_u16_u16_205_wire;
    -- flow-through select operator MUX_208_inst
    n_winr_209 <= MUX_206_wire when (flag1_188(0) /=  '0') else winr_66;
    -- flow-through select operator MUX_219_inst
    MUX_219_wire <= konst_215_wire_constant when (col_done_198(0) /=  '0') else ADD_u16_u16_218_wire;
    -- flow-through select operator MUX_221_inst
    n_col_222 <= MUX_219_wire when (AND_u1_u1_213_wire(0) /=  '0') else col_71;
    -- flow-through select operator MUX_233_inst
    n_row_234 <= ADD_u16_u16_231_wire when (AND_u1_u1_228_wire(0) /=  '0') else row_76;
    -- flow-through select operator MUX_268_inst
    n_word_start_269 <= type_cast_266_wire when (flag1_188(0) /=  '0') else konst_267_wire_constant;
    -- flow-through select operator MUX_279_inst
    n_address_280 <= type_cast_275_wire when (flag1_188(0) /=  '0') else ADD_u64_u64_278_wire;
    -- flow-through select operator MUX_287_inst
    n_left_288 <= nl_start_35 when (flag1_188(0) /=  '0') else SUB_u16_u16_286_wire;
    -- flow-through select operator MUX_300_inst
    MUX_300_wire <= SUB_u16_u16_298_wire when (UGT_u16_u1_295_wire(0) /=  '0') else fn_blk_43;
    -- flow-through select operator MUX_306_inst
    MUX_306_wire <= n_left_288 when (ULT_u16_u1_303_wire(0) /=  '0') else konst_305_wire_constant;
    -- flow-through select operator MUX_307_inst
    n_blk_308 <= MUX_300_wire when (flag1_188(0) /=  '0') else MUX_306_wire;
    -- flow-through select operator MUX_42_inst
    fn_blk_43 <= num_cont_buffer when (ULT_u16_u1_39_wire(0) /=  '0') else konst_41_wire_constant;
    slice_142_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_142_inst_req_0;
      slice_142_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_142_inst_req_1;
      slice_142_inst_ack_1<= update_ack(0);
      slice_142_inst: SliceSplitProtocol generic map(name => "slice_142_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w1_143, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_146_inst_req_0;
      slice_146_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_146_inst_req_1;
      slice_146_inst_ack_1<= update_ack(0);
      slice_146_inst: SliceSplitProtocol generic map(name => "slice_146_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w2_147, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_150_inst_req_0;
      slice_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_150_inst_req_1;
      slice_150_inst_ack_1<= update_ack(0);
      slice_150_inst: SliceSplitProtocol generic map(name => "slice_150_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w3_151, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_154_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_154_inst_req_0;
      slice_154_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_154_inst_req_1;
      slice_154_inst_ack_1<= update_ack(0);
      slice_154_inst: SliceSplitProtocol generic map(name => "slice_154_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w4_155, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_156_delayed_14_0_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_156_delayed_14_0_156_inst_req_0;
      W_c1_156_delayed_14_0_156_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_156_delayed_14_0_156_inst_req_1;
      W_c1_156_delayed_14_0_156_inst_ack_1<= rack(0);
      W_c1_156_delayed_14_0_156_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_156_delayed_14_0_156_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_156_delayed_14_0_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_160_delayed_14_0_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_160_delayed_14_0_163_inst_req_0;
      W_c2_160_delayed_14_0_163_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_160_delayed_14_0_163_inst_req_1;
      W_c2_160_delayed_14_0_163_inst_ack_1<= rack(0);
      W_c2_160_delayed_14_0_163_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_160_delayed_14_0_163_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_160_delayed_14_0_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_164_delayed_14_0_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_164_delayed_14_0_170_inst_req_0;
      W_c3_164_delayed_14_0_170_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_164_delayed_14_0_170_inst_req_1;
      W_c3_164_delayed_14_0_170_inst_ack_1<= rack(0);
      W_c3_164_delayed_14_0_170_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_164_delayed_14_0_170_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_164_delayed_14_0_172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_168_delayed_14_0_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_168_delayed_14_0_177_inst_req_0;
      W_c4_168_delayed_14_0_177_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_168_delayed_14_0_177_inst_req_1;
      W_c4_168_delayed_14_0_177_inst_ack_1<= rack(0);
      W_c4_168_delayed_14_0_177_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_168_delayed_14_0_177_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_168_delayed_14_0_179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_33_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_35 <= tmp_var; -- 
    end process;
    addr_of_134_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_134_final_reg_req_0;
      addr_of_134_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_134_final_reg_req_1;
      addr_of_134_final_reg_ack_1<= rack(0);
      addr_of_134_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_134_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_133_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_280_50_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_280_50_buf_req_0;
      n_address_280_50_buf_ack_0<= wack(0);
      rreq(0) <= n_address_280_50_buf_req_1;
      n_address_280_50_buf_ack_1<= rack(0);
      n_address_280_50_buf : InterlockBuffer generic map ( -- 
        name => "n_address_280_50_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_280_50_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_308_65_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_308_65_buf_req_0;
      n_blk_308_65_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_308_65_buf_req_1;
      n_blk_308_65_buf_ack_1<= rack(0);
      n_blk_308_65_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_308_65_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_308_65_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_222_75_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_222_75_buf_req_0;
      n_col_222_75_buf_ack_0<= wack(0);
      rreq(0) <= n_col_222_75_buf_req_1;
      n_col_222_75_buf_ack_1<= rack(0);
      n_col_222_75_buf : InterlockBuffer generic map ( -- 
        name => "n_col_222_75_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_222_75_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_288_60_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_288_60_buf_req_0;
      n_left_288_60_buf_ack_0<= wack(0);
      rreq(0) <= n_left_288_60_buf_req_1;
      n_left_288_60_buf_ack_1<= rack(0);
      n_left_288_60_buf : InterlockBuffer generic map ( -- 
        name => "n_left_288_60_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_288_60_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_234_78_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_234_78_buf_req_0;
      n_row_234_78_buf_ack_0<= wack(0);
      rreq(0) <= n_row_234_78_buf_req_1;
      n_row_234_78_buf_ack_1<= rack(0);
      n_row_234_78_buf : InterlockBuffer generic map ( -- 
        name => "n_row_234_78_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_234_78_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_209_70_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_209_70_buf_req_0;
      n_winr_209_70_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_209_70_buf_req_1;
      n_winr_209_70_buf_ack_1<= rack(0);
      n_winr_209_70_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_209_70_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_209_70_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_269_56_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_269_56_buf_req_0;
      n_word_start_269_56_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_269_56_buf_req_1;
      n_word_start_269_56_buf_ack_1<= rack(0);
      n_word_start_269_56_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_269_56_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_269_56_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_35_59_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_35_59_buf_req_0;
      nl_start_35_59_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_35_59_buf_req_1;
      nl_start_35_59_buf_ack_1<= rack(0);
      nl_start_35_59_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_35_59_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_35_59_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_124_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_51(1 downto 0);
      type_cast_124_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_243_inst
    process(MUL_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_242_wire(15 downto 0);
      na1_244 <= tmp_var; -- 
    end process;
    -- interlock type_cast_248_inst
    process(n_winr_209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_209(15 downto 0);
      type_cast_248_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_250_inst
    process(MUL_u32_u32_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_249_wire(31 downto 0);
      na2_251 <= tmp_var; -- 
    end process;
    -- interlock type_cast_261_inst
    process(AND_u32_u32_260_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_260_wire(15 downto 0);
      na4_262 <= tmp_var; -- 
    end process;
    -- interlock type_cast_266_inst
    process(na4_262) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_262(1 downto 0);
      type_cast_266_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_275_inst
    process(LSHR_u32_u32_274_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_274_wire(31 downto 0);
      type_cast_275_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_31_inst
    process(MUL_u16_u16_30_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_30_wire(15 downto 0);
      m_factor_32 <= tmp_var; -- 
    end process;
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_43,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_64_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_133_index_1_rename
    process(R_address_132_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_132_resized;
      ov(13 downto 0) := iv;
      R_address_132_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_index_1_resize
    process(address_46) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_46;
      ov := iv(13 downto 0);
      R_address_132_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_root_address_inst
    process(array_obj_ref_133_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_133_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_addr_0
    process(ptr_deref_138_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_base_resize
    process(fetch_addr_135) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_135;
      ov := iv(13 downto 0);
      ptr_deref_138_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_gather_scatter
    process(ptr_deref_138_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_data_0;
      ov(63 downto 0) := iv;
      word_read_139 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_root_address_inst
    process(ptr_deref_138_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_44_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_312_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_44_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_44_branch_req_0,
          ack0 => do_while_stmt_44_branch_ack_0,
          ack1 => do_while_stmt_44_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_125_inst
    process(num_blk_61, type_cast_124_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_61, type_cast_124_wire, tmp_var);
      ADD_u16_u16_125_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_205_inst
    process(winr_66) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_66, konst_204_wire_constant, tmp_var);
      ADD_u16_u16_205_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_218_inst
    process(col_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_71, konst_217_wire_constant, tmp_var);
      ADD_u16_u16_218_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_231_inst
    process(row_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_76, konst_230_wire_constant, tmp_var);
      ADD_u16_u16_231_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_241_inst
    process(n_col_222, MUL_u16_u16_240_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_222, MUL_u16_u16_240_wire, tmp_var);
      ADD_u16_u16_241_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_293_inst
    process(fn_blk_43, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_43, na4_262, tmp_var);
      ADD_u16_u16_293_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_255_inst
    process(na1_244, na2_251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_244, na2_251, tmp_var);
      na3_256 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_278_inst
    process(address_46) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_46, konst_277_wire_constant, tmp_var);
      ADD_u64_u64_278_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_107_inst
    process(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire, tmp_var);
      AND_u1_u1_107_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_114_inst
    process(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire, tmp_var);
      AND_u1_u1_114_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_213_inst
    process(winr_done_193, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, flag1_188, tmp_var);
      AND_u1_u1_213_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_227_inst
    process(col_done_198, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_198, flag1_188, tmp_var);
      AND_u1_u1_227_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_228_inst
    process(winr_done_193, AND_u1_u1_227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, AND_u1_u1_227_wire, tmp_var);
      AND_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_94_inst
    process(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire, tmp_var);
      AND_u1_u1_94_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_260_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_256, konst_259_wire_constant, tmp_var);
      AND_u32_u32_260_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_187_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_57, num_blk_61, tmp_var);
      flag1_188 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_192_inst
    process(winr_66, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_66, rk1_buffer, tmp_var);
      winr_done_193 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_197_inst
    process(col_71, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_71, col1_buffer, tmp_var);
      col_done_198 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_103_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_102_wire_constant, tmp_var);
      EQ_u2_u1_103_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_110_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_109_wire_constant, tmp_var);
      EQ_u2_u1_110_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_117_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_116_wire_constant, tmp_var);
      EQ_u2_u1_117_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_85_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_84_wire_constant, tmp_var);
      c1_86 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_90_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_89_wire_constant, tmp_var);
      EQ_u2_u1_90_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_97_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_96_wire_constant, tmp_var);
      EQ_u2_u1_97_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_274_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_256, konst_273_wire_constant, tmp_var);
      LSHR_u32_u32_274_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_240_inst
    process(ct_buffer, n_row_234) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_234, tmp_var);
      MUL_u16_u16_240_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_242_inst
    process(chl_in_buffer, ADD_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_241_wire, tmp_var);
      MUL_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_30_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_30_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(m_factor_32, type_cast_248_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_32, type_cast_248_wire, tmp_var);
      MUL_u32_u32_249_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_312_inst
    process(n_row_234, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_234, row1_buffer, tmp_var);
      NEQ_u16_u1_312_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_118_inst
    process(AND_u1_u1_114_wire, EQ_u2_u1_117_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_114_wire, EQ_u2_u1_117_wire, tmp_var);
      OR_u1_u1_118_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_119_inst
    process(AND_u1_u1_107_wire, OR_u1_u1_118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_107_wire, OR_u1_u1_118_wire, tmp_var);
      c3_120 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_98_inst
    process(AND_u1_u1_94_wire, EQ_u2_u1_97_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_94_wire, EQ_u2_u1_97_wire, tmp_var);
      c2_99 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_286_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_57, num_blk_61, tmp_var);
      SUB_u16_u16_286_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_298_inst
    process(konst_296_wire_constant, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_296_wire_constant, na4_262, tmp_var);
      SUB_u16_u16_298_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_106_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_105_wire_constant, tmp_var);
      UGT_u16_u1_106_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_113_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_112_wire_constant, tmp_var);
      UGT_u16_u1_113_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_127_inst
    process(ADD_u16_u16_125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_125_wire, konst_126_wire_constant, tmp_var);
      c4_128 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_295_inst
    process(ADD_u16_u16_293_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_293_wire, konst_294_wire_constant, tmp_var);
      UGT_u16_u1_295_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_93_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_92_wire_constant, tmp_var);
      UGT_u16_u1_93_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_303_inst
    process(n_left_288) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_288, konst_302_wire_constant, tmp_var);
      ULT_u16_u1_303_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_39_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_38_wire_constant, tmp_var);
      ULT_u16_u1_39_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_133_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_132_scaled;
      array_obj_ref_133_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_133_index_offset_req_0;
      array_obj_ref_133_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_133_index_offset_req_1;
      array_obj_ref_133_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_138_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_138_load_0_req_0;
      ptr_deref_138_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_138_load_0_req_1;
      ptr_deref_138_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_138_word_address_0;
      ptr_deref_138_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_167_inst WPIPE_input_pipe1_160_inst WPIPE_input_pipe1_174_inst WPIPE_input_pipe1_181_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_167_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_160_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_174_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_0;
      WPIPE_input_pipe1_167_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_160_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_174_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_167_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_160_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_174_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_1;
      WPIPE_input_pipe1_167_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_160_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_174_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_168_delayed_14_0_179(0);
      guard_vector(1)  <= c3_164_delayed_14_0_172(0);
      guard_vector(2)  <= c1_156_delayed_14_0_158(0);
      guard_vector(3)  <= c2_160_delayed_14_0_165(0);
      data_in <= w2_147 & w1_143 & w3_151 & w4_155;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1120_start: Boolean;
  signal convolution3D_CP_1120_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_518_inst_ack_0 : boolean;
  signal type_cast_543_inst_req_0 : boolean;
  signal type_cast_660_inst_ack_0 : boolean;
  signal type_cast_506_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_502_inst_ack_1 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_564_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_589_inst_ack_1 : boolean;
  signal type_cast_568_inst_ack_1 : boolean;
  signal type_cast_506_inst_ack_0 : boolean;
  signal type_cast_618_inst_req_0 : boolean;
  signal type_cast_606_inst_req_1 : boolean;
  signal type_cast_631_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_502_inst_ack_0 : boolean;
  signal type_cast_606_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_589_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_527_inst_ack_0 : boolean;
  signal type_cast_568_inst_ack_0 : boolean;
  signal type_cast_531_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_589_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_564_inst_req_1 : boolean;
  signal type_cast_581_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_577_inst_req_1 : boolean;
  signal type_cast_631_inst_ack_0 : boolean;
  signal type_cast_618_inst_ack_1 : boolean;
  signal type_cast_640_inst_req_1 : boolean;
  signal type_cast_518_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_552_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_req_0 : boolean;
  signal type_cast_660_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_577_inst_ack_1 : boolean;
  signal type_cast_543_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_552_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_502_inst_req_0 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_502_inst_req_1 : boolean;
  signal type_cast_631_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_514_inst_ack_1 : boolean;
  signal type_cast_618_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_589_inst_req_0 : boolean;
  signal type_cast_568_inst_req_1 : boolean;
  signal type_cast_568_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_602_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_602_inst_ack_0 : boolean;
  signal type_cast_531_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_552_inst_ack_0 : boolean;
  signal type_cast_644_inst_req_0 : boolean;
  signal type_cast_644_inst_req_1 : boolean;
  signal type_cast_640_inst_ack_1 : boolean;
  signal type_cast_644_inst_ack_1 : boolean;
  signal type_cast_618_inst_ack_0 : boolean;
  signal type_cast_543_inst_ack_1 : boolean;
  signal type_cast_606_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_527_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_614_inst_ack_1 : boolean;
  signal type_cast_644_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_577_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_552_inst_req_0 : boolean;
  signal type_cast_631_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_ack_0 : boolean;
  signal type_cast_543_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_527_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_527_inst_ack_1 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal type_cast_556_inst_req_0 : boolean;
  signal type_cast_606_inst_ack_1 : boolean;
  signal type_cast_506_inst_req_1 : boolean;
  signal type_cast_556_inst_ack_0 : boolean;
  signal type_cast_581_inst_req_1 : boolean;
  signal addr_of_1228_final_reg_req_1 : boolean;
  signal type_cast_556_inst_req_1 : boolean;
  signal type_cast_556_inst_ack_1 : boolean;
  signal type_cast_640_inst_req_0 : boolean;
  signal type_cast_531_inst_req_0 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal type_cast_506_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_614_inst_req_0 : boolean;
  signal type_cast_1338_inst_ack_0 : boolean;
  signal type_cast_688_inst_req_0 : boolean;
  signal type_cast_688_inst_ack_0 : boolean;
  signal addr_of_1228_final_reg_ack_0 : boolean;
  signal addr_of_1228_final_reg_req_0 : boolean;
  signal type_cast_1338_inst_req_0 : boolean;
  signal type_cast_1248_inst_req_1 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal type_cast_581_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_627_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_577_inst_req_0 : boolean;
  signal type_cast_1302_inst_req_1 : boolean;
  signal type_cast_688_inst_req_1 : boolean;
  signal type_cast_688_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_627_inst_req_1 : boolean;
  signal type_cast_1248_inst_ack_0 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_713_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_ack_1 : boolean;
  signal type_cast_713_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_564_inst_ack_0 : boolean;
  signal type_cast_704_inst_req_0 : boolean;
  signal type_cast_704_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_514_inst_req_1 : boolean;
  signal type_cast_660_inst_ack_1 : boolean;
  signal type_cast_1248_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_req_1 : boolean;
  signal type_cast_660_inst_req_1 : boolean;
  signal if_stmt_668_branch_ack_0 : boolean;
  signal if_stmt_668_branch_ack_1 : boolean;
  signal if_stmt_668_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_514_inst_ack_0 : boolean;
  signal type_cast_704_inst_req_1 : boolean;
  signal type_cast_704_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_614_inst_req_1 : boolean;
  signal type_cast_581_inst_req_0 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal type_cast_713_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_req_1 : boolean;
  signal type_cast_713_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1231_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_602_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_627_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_514_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_564_inst_req_0 : boolean;
  signal addr_of_1228_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_627_inst_req_0 : boolean;
  signal type_cast_518_inst_ack_1 : boolean;
  signal type_cast_640_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_539_inst_req_1 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal type_cast_531_inst_ack_0 : boolean;
  signal type_cast_518_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1231_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_602_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1231_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1231_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_439_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_439_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_439_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_439_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_req_0 : boolean;
  signal type_cast_443_inst_req_0 : boolean;
  signal type_cast_443_inst_ack_0 : boolean;
  signal type_cast_443_inst_req_1 : boolean;
  signal type_cast_443_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_req_0 : boolean;
  signal type_cast_1284_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_req_1 : boolean;
  signal type_cast_1284_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_452_inst_ack_1 : boolean;
  signal type_cast_456_inst_req_0 : boolean;
  signal type_cast_456_inst_ack_0 : boolean;
  signal type_cast_456_inst_req_1 : boolean;
  signal type_cast_456_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_464_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_464_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_464_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_464_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_614_inst_ack_0 : boolean;
  signal type_cast_468_inst_req_0 : boolean;
  signal type_cast_468_inst_ack_0 : boolean;
  signal type_cast_468_inst_req_1 : boolean;
  signal type_cast_468_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_477_inst_ack_1 : boolean;
  signal type_cast_481_inst_req_0 : boolean;
  signal type_cast_481_inst_ack_0 : boolean;
  signal type_cast_481_inst_req_1 : boolean;
  signal type_cast_481_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_489_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_489_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_489_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_489_inst_ack_1 : boolean;
  signal type_cast_493_inst_req_0 : boolean;
  signal type_cast_493_inst_ack_0 : boolean;
  signal type_cast_493_inst_req_1 : boolean;
  signal type_cast_493_inst_ack_1 : boolean;
  signal type_cast_1248_inst_req_0 : boolean;
  signal type_cast_723_inst_req_0 : boolean;
  signal type_cast_723_inst_ack_0 : boolean;
  signal type_cast_723_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_ack_0 : boolean;
  signal type_cast_723_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_req_0 : boolean;
  signal type_cast_1302_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1244_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1244_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1244_inst_ack_0 : boolean;
  signal type_cast_1302_inst_ack_0 : boolean;
  signal array_obj_ref_758_index_offset_req_0 : boolean;
  signal array_obj_ref_758_index_offset_ack_0 : boolean;
  signal array_obj_ref_758_index_offset_req_1 : boolean;
  signal array_obj_ref_758_index_offset_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1244_inst_req_0 : boolean;
  signal array_obj_ref_1227_index_offset_ack_1 : boolean;
  signal addr_of_759_final_reg_req_0 : boolean;
  signal addr_of_759_final_reg_ack_0 : boolean;
  signal addr_of_759_final_reg_req_1 : boolean;
  signal addr_of_759_final_reg_ack_1 : boolean;
  signal array_obj_ref_1227_index_offset_req_1 : boolean;
  signal type_cast_1302_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_762_inst_req_0 : boolean;
  signal type_cast_1266_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_762_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_762_inst_req_1 : boolean;
  signal type_cast_1266_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_762_inst_ack_1 : boolean;
  signal type_cast_1338_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_req_0 : boolean;
  signal type_cast_766_inst_req_0 : boolean;
  signal type_cast_766_inst_ack_0 : boolean;
  signal type_cast_766_inst_req_1 : boolean;
  signal type_cast_766_inst_ack_1 : boolean;
  signal array_obj_ref_1227_index_offset_ack_0 : boolean;
  signal type_cast_1284_inst_ack_1 : boolean;
  signal array_obj_ref_1227_index_offset_req_0 : boolean;
  signal type_cast_1284_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_775_inst_req_0 : boolean;
  signal type_cast_1266_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_775_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_775_inst_req_1 : boolean;
  signal type_cast_1266_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_775_inst_ack_1 : boolean;
  signal type_cast_1235_inst_ack_1 : boolean;
  signal type_cast_1235_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_ack_1 : boolean;
  signal type_cast_779_inst_req_0 : boolean;
  signal type_cast_779_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_req_1 : boolean;
  signal type_cast_779_inst_req_1 : boolean;
  signal type_cast_779_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_ack_1 : boolean;
  signal type_cast_1235_inst_ack_0 : boolean;
  signal type_cast_1235_inst_req_0 : boolean;
  signal type_cast_797_inst_req_0 : boolean;
  signal type_cast_797_inst_ack_0 : boolean;
  signal type_cast_797_inst_req_1 : boolean;
  signal type_cast_797_inst_ack_1 : boolean;
  signal type_cast_1460_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_ack_1 : boolean;
  signal type_cast_815_inst_req_0 : boolean;
  signal type_cast_815_inst_ack_0 : boolean;
  signal type_cast_815_inst_req_1 : boolean;
  signal type_cast_752_inst_req_0 : boolean;
  signal type_cast_815_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_ack_0 : boolean;
  signal type_cast_1518_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_ack_1 : boolean;
  signal type_cast_833_inst_req_0 : boolean;
  signal type_cast_833_inst_ack_0 : boolean;
  signal type_cast_833_inst_req_1 : boolean;
  signal type_cast_833_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_ack_1 : boolean;
  signal type_cast_994_inst_req_0 : boolean;
  signal type_cast_994_inst_ack_0 : boolean;
  signal type_cast_1467_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_ack_1 : boolean;
  signal type_cast_943_inst_req_0 : boolean;
  signal type_cast_1518_inst_req_1 : boolean;
  signal type_cast_943_inst_ack_0 : boolean;
  signal type_cast_869_inst_req_0 : boolean;
  signal type_cast_869_inst_ack_0 : boolean;
  signal type_cast_869_inst_req_1 : boolean;
  signal type_cast_869_inst_ack_1 : boolean;
  signal type_cast_1221_inst_req_0 : boolean;
  signal phi_stmt_1454_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_ack_1 : boolean;
  signal type_cast_1467_inst_req_1 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal type_cast_1221_inst_ack_0 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal type_cast_943_inst_req_1 : boolean;
  signal phi_stmt_1409_req_1 : boolean;
  signal type_cast_943_inst_ack_1 : boolean;
  signal phi_stmt_1409_ack_0 : boolean;
  signal type_cast_994_inst_req_1 : boolean;
  signal type_cast_752_inst_ack_0 : boolean;
  signal type_cast_994_inst_ack_1 : boolean;
  signal type_cast_1221_inst_req_1 : boolean;
  signal type_cast_1467_inst_ack_1 : boolean;
  signal phi_stmt_988_req_1 : boolean;
  signal ptr_deref_895_store_0_req_0 : boolean;
  signal ptr_deref_895_store_0_ack_0 : boolean;
  signal ptr_deref_895_store_0_req_1 : boolean;
  signal ptr_deref_895_store_0_ack_1 : boolean;
  signal phi_stmt_940_req_0 : boolean;
  signal phi_stmt_981_ack_0 : boolean;
  signal phi_stmt_988_ack_0 : boolean;
  signal type_cast_752_inst_req_1 : boolean;
  signal if_stmt_909_branch_req_0 : boolean;
  signal type_cast_752_inst_ack_1 : boolean;
  signal if_stmt_909_branch_ack_1 : boolean;
  signal if_stmt_909_branch_ack_0 : boolean;
  signal phi_stmt_746_req_1 : boolean;
  signal phi_stmt_1461_req_1 : boolean;
  signal if_stmt_960_branch_req_0 : boolean;
  signal if_stmt_960_branch_ack_1 : boolean;
  signal if_stmt_960_branch_ack_0 : boolean;
  signal type_cast_1518_inst_ack_1 : boolean;
  signal type_cast_1221_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1009_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1009_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1009_inst_req_1 : boolean;
  signal phi_stmt_1215_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1009_inst_ack_1 : boolean;
  signal phi_stmt_1515_req_0 : boolean;
  signal phi_stmt_940_ack_0 : boolean;
  signal type_cast_1013_inst_req_0 : boolean;
  signal type_cast_1013_inst_ack_0 : boolean;
  signal type_cast_1013_inst_req_1 : boolean;
  signal type_cast_1013_inst_ack_1 : boolean;
  signal phi_stmt_746_ack_0 : boolean;
  signal type_cast_1028_inst_req_0 : boolean;
  signal type_cast_1028_inst_ack_0 : boolean;
  signal type_cast_1028_inst_req_1 : boolean;
  signal type_cast_1028_inst_ack_1 : boolean;
  signal phi_stmt_1461_req_0 : boolean;
  signal if_stmt_1035_branch_req_0 : boolean;
  signal if_stmt_1035_branch_ack_1 : boolean;
  signal if_stmt_1035_branch_ack_0 : boolean;
  signal array_obj_ref_1074_index_offset_req_0 : boolean;
  signal array_obj_ref_1074_index_offset_ack_0 : boolean;
  signal array_obj_ref_1074_index_offset_req_1 : boolean;
  signal array_obj_ref_1074_index_offset_ack_1 : boolean;
  signal addr_of_1075_final_reg_req_0 : boolean;
  signal addr_of_1075_final_reg_ack_0 : boolean;
  signal addr_of_1075_final_reg_req_1 : boolean;
  signal addr_of_1075_final_reg_ack_1 : boolean;
  signal ptr_deref_1078_store_0_req_0 : boolean;
  signal ptr_deref_1078_store_0_ack_0 : boolean;
  signal ptr_deref_1078_store_0_req_1 : boolean;
  signal ptr_deref_1078_store_0_ack_1 : boolean;
  signal type_cast_1085_inst_req_0 : boolean;
  signal type_cast_1085_inst_ack_0 : boolean;
  signal type_cast_1085_inst_req_1 : boolean;
  signal type_cast_1085_inst_ack_1 : boolean;
  signal type_cast_1089_inst_req_0 : boolean;
  signal type_cast_1089_inst_ack_0 : boolean;
  signal type_cast_1089_inst_req_1 : boolean;
  signal type_cast_1089_inst_ack_1 : boolean;
  signal type_cast_1093_inst_req_0 : boolean;
  signal type_cast_1093_inst_ack_0 : boolean;
  signal type_cast_1093_inst_req_1 : boolean;
  signal type_cast_1093_inst_ack_1 : boolean;
  signal type_cast_1097_inst_req_0 : boolean;
  signal type_cast_1097_inst_ack_0 : boolean;
  signal type_cast_1097_inst_req_1 : boolean;
  signal type_cast_1097_inst_ack_1 : boolean;
  signal if_stmt_1135_branch_req_0 : boolean;
  signal if_stmt_1135_branch_ack_1 : boolean;
  signal if_stmt_1135_branch_ack_0 : boolean;
  signal type_cast_1156_inst_req_0 : boolean;
  signal type_cast_1156_inst_ack_0 : boolean;
  signal type_cast_1156_inst_req_1 : boolean;
  signal type_cast_1156_inst_ack_1 : boolean;
  signal type_cast_1160_inst_req_0 : boolean;
  signal type_cast_1160_inst_ack_0 : boolean;
  signal type_cast_1160_inst_req_1 : boolean;
  signal type_cast_1160_inst_ack_1 : boolean;
  signal type_cast_1169_inst_req_0 : boolean;
  signal type_cast_1169_inst_ack_0 : boolean;
  signal type_cast_1169_inst_req_1 : boolean;
  signal type_cast_1169_inst_ack_1 : boolean;
  signal type_cast_1178_inst_req_0 : boolean;
  signal type_cast_1178_inst_ack_0 : boolean;
  signal type_cast_1178_inst_req_1 : boolean;
  signal type_cast_1178_inst_ack_1 : boolean;
  signal type_cast_1187_inst_req_0 : boolean;
  signal type_cast_1187_inst_ack_0 : boolean;
  signal type_cast_1187_inst_req_1 : boolean;
  signal type_cast_1187_inst_ack_1 : boolean;
  signal type_cast_1192_inst_req_0 : boolean;
  signal type_cast_1192_inst_ack_0 : boolean;
  signal type_cast_1192_inst_req_1 : boolean;
  signal type_cast_1192_inst_ack_1 : boolean;
  signal type_cast_1338_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_ack_1 : boolean;
  signal type_cast_1356_inst_req_0 : boolean;
  signal type_cast_1356_inst_ack_0 : boolean;
  signal type_cast_1356_inst_req_1 : boolean;
  signal type_cast_1356_inst_ack_1 : boolean;
  signal ptr_deref_1364_store_0_req_0 : boolean;
  signal ptr_deref_1364_store_0_ack_0 : boolean;
  signal ptr_deref_1364_store_0_req_1 : boolean;
  signal ptr_deref_1364_store_0_ack_1 : boolean;
  signal if_stmt_1378_branch_req_0 : boolean;
  signal if_stmt_1378_branch_ack_1 : boolean;
  signal if_stmt_1378_branch_ack_0 : boolean;
  signal if_stmt_1429_branch_req_0 : boolean;
  signal if_stmt_1429_branch_ack_1 : boolean;
  signal if_stmt_1429_branch_ack_0 : boolean;
  signal type_cast_1045_inst_ack_0 : boolean;
  signal type_cast_1045_inst_req_0 : boolean;
  signal type_cast_1467_inst_req_0 : boolean;
  signal type_cast_1444_inst_req_0 : boolean;
  signal type_cast_1444_inst_ack_0 : boolean;
  signal type_cast_1444_inst_req_1 : boolean;
  signal type_cast_1444_inst_ack_1 : boolean;
  signal type_cast_1518_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1482_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1482_inst_ack_0 : boolean;
  signal phi_stmt_1409_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1482_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1482_inst_ack_1 : boolean;
  signal type_cast_1412_inst_ack_1 : boolean;
  signal phi_stmt_981_req_1 : boolean;
  signal type_cast_1486_inst_req_0 : boolean;
  signal type_cast_1486_inst_ack_0 : boolean;
  signal type_cast_1486_inst_req_1 : boolean;
  signal type_cast_1486_inst_ack_1 : boolean;
  signal type_cast_1412_inst_req_1 : boolean;
  signal type_cast_987_inst_ack_1 : boolean;
  signal type_cast_1501_inst_req_0 : boolean;
  signal type_cast_1501_inst_ack_0 : boolean;
  signal type_cast_1501_inst_req_1 : boolean;
  signal phi_stmt_1215_req_0 : boolean;
  signal type_cast_1501_inst_ack_1 : boolean;
  signal type_cast_987_inst_req_1 : boolean;
  signal if_stmt_1508_branch_req_0 : boolean;
  signal if_stmt_1508_branch_ack_1 : boolean;
  signal if_stmt_1508_branch_ack_0 : boolean;
  signal type_cast_1412_inst_ack_0 : boolean;
  signal type_cast_1412_inst_req_0 : boolean;
  signal type_cast_987_inst_ack_0 : boolean;
  signal type_cast_987_inst_req_0 : boolean;
  signal array_obj_ref_1547_index_offset_req_0 : boolean;
  signal array_obj_ref_1547_index_offset_ack_0 : boolean;
  signal array_obj_ref_1547_index_offset_req_1 : boolean;
  signal array_obj_ref_1547_index_offset_ack_1 : boolean;
  signal addr_of_1548_final_reg_req_0 : boolean;
  signal addr_of_1548_final_reg_ack_0 : boolean;
  signal addr_of_1548_final_reg_req_1 : boolean;
  signal addr_of_1548_final_reg_ack_1 : boolean;
  signal ptr_deref_1551_store_0_req_0 : boolean;
  signal ptr_deref_1551_store_0_ack_0 : boolean;
  signal ptr_deref_1551_store_0_req_1 : boolean;
  signal ptr_deref_1551_store_0_ack_1 : boolean;
  signal phi_stmt_1515_ack_0 : boolean;
  signal call_stmt_1558_call_req_0 : boolean;
  signal call_stmt_1558_call_ack_0 : boolean;
  signal call_stmt_1558_call_req_1 : boolean;
  signal call_stmt_1558_call_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1570_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1570_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1570_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1570_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1573_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1573_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1573_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1573_inst_ack_1 : boolean;
  signal phi_stmt_988_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1577_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1577_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1577_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1577_inst_ack_1 : boolean;
  signal phi_stmt_1461_ack_0 : boolean;
  signal phi_stmt_1454_ack_0 : boolean;
  signal phi_stmt_981_req_0 : boolean;
  signal phi_stmt_1454_req_1 : boolean;
  signal type_cast_1601_inst_req_0 : boolean;
  signal phi_stmt_1042_ack_0 : boolean;
  signal type_cast_1601_inst_ack_0 : boolean;
  signal type_cast_1460_inst_ack_1 : boolean;
  signal type_cast_1601_inst_req_1 : boolean;
  signal type_cast_1601_inst_ack_1 : boolean;
  signal phi_stmt_940_req_1 : boolean;
  signal type_cast_1460_inst_req_1 : boolean;
  signal type_cast_1611_inst_req_0 : boolean;
  signal type_cast_1611_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_1 : boolean;
  signal phi_stmt_1042_req_0 : boolean;
  signal type_cast_1611_inst_ack_1 : boolean;
  signal phi_stmt_1215_ack_0 : boolean;
  signal type_cast_1620_inst_req_0 : boolean;
  signal type_cast_1045_inst_ack_1 : boolean;
  signal type_cast_1620_inst_ack_0 : boolean;
  signal type_cast_1460_inst_ack_0 : boolean;
  signal type_cast_1620_inst_req_1 : boolean;
  signal type_cast_1045_inst_req_1 : boolean;
  signal type_cast_1620_inst_ack_1 : boolean;
  signal type_cast_1649_inst_req_0 : boolean;
  signal type_cast_1649_inst_ack_0 : boolean;
  signal type_cast_1649_inst_req_1 : boolean;
  signal type_cast_1649_inst_ack_1 : boolean;
  signal type_cast_1653_inst_req_0 : boolean;
  signal type_cast_1653_inst_ack_0 : boolean;
  signal type_cast_1653_inst_req_1 : boolean;
  signal type_cast_1653_inst_ack_1 : boolean;
  signal call_stmt_1657_call_req_0 : boolean;
  signal call_stmt_1657_call_ack_0 : boolean;
  signal call_stmt_1657_call_req_1 : boolean;
  signal call_stmt_1657_call_ack_1 : boolean;
  signal call_stmt_1664_call_req_0 : boolean;
  signal call_stmt_1664_call_ack_0 : boolean;
  signal call_stmt_1664_call_req_1 : boolean;
  signal call_stmt_1664_call_ack_1 : boolean;
  signal if_stmt_1676_branch_req_0 : boolean;
  signal if_stmt_1676_branch_ack_1 : boolean;
  signal if_stmt_1676_branch_ack_0 : boolean;
  signal type_cast_1686_inst_req_0 : boolean;
  signal type_cast_1686_inst_ack_0 : boolean;
  signal type_cast_1686_inst_req_1 : boolean;
  signal type_cast_1686_inst_ack_1 : boolean;
  signal call_stmt_1690_call_req_0 : boolean;
  signal call_stmt_1690_call_ack_0 : boolean;
  signal call_stmt_1690_call_req_1 : boolean;
  signal call_stmt_1690_call_ack_1 : boolean;
  signal type_cast_1694_inst_req_0 : boolean;
  signal type_cast_1694_inst_ack_0 : boolean;
  signal type_cast_1694_inst_req_1 : boolean;
  signal type_cast_1694_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1701_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1701_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1701_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1701_inst_ack_1 : boolean;
  signal phi_stmt_746_req_0 : boolean;
  signal phi_stmt_1629_req_1 : boolean;
  signal type_cast_1632_inst_req_0 : boolean;
  signal type_cast_1632_inst_ack_0 : boolean;
  signal type_cast_1632_inst_req_1 : boolean;
  signal type_cast_1632_inst_ack_1 : boolean;
  signal phi_stmt_1629_req_0 : boolean;
  signal phi_stmt_1629_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1120_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1120: Block -- control-path 
    signal convolution3D_CP_1120_elements: BooleanArray(335 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1120_elements(0) <= convolution3D_CP_1120_start;
    convolution3D_CP_1120_symbol <= convolution3D_CP_1120_elements(267);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_436/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/branch_block_stmt_436__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Update/cr
      -- 
    cr_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_606_inst_req_1); -- 
    cr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_640_inst_req_1); -- 
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_543_inst_req_1); -- 
    cr_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_593_inst_req_1); -- 
    cr_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_618_inst_req_1); -- 
    cr_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_568_inst_req_1); -- 
    cr_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_531_inst_req_1); -- 
    cr_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_644_inst_req_1); -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_631_inst_req_1); -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_506_inst_req_1); -- 
    cr_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_581_inst_req_1); -- 
    cr_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_556_inst_req_1); -- 
    cr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_660_inst_req_1); -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_518_inst_req_1); -- 
    rr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => RPIPE_maxpool_input_pipe_439_inst_req_0); -- 
    cr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_443_inst_req_1); -- 
    cr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_456_inst_req_1); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_468_inst_req_1); -- 
    cr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_481_inst_req_1); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_493_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_update_start_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Update/cr
      -- 
    ra_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_439_inst_ack_0, ack => convolution3D_CP_1120_elements(1)); -- 
    cr_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(1), ack => RPIPE_maxpool_input_pipe_439_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_439_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Sample/rr
      -- 
    ca_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_439_inst_ack_1, ack => convolution3D_CP_1120_elements(2)); -- 
    rr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => type_cast_443_inst_req_0); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => RPIPE_maxpool_input_pipe_452_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Sample/ra
      -- 
    ra_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_0, ack => convolution3D_CP_1120_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_443_Update/ca
      -- 
    ca_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_1, ack => convolution3D_CP_1120_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_update_start_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Update/cr
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_452_inst_ack_0, ack => convolution3D_CP_1120_elements(5)); -- 
    cr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(5), ack => RPIPE_maxpool_input_pipe_452_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_452_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Sample/rr
      -- 
    ca_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_452_inst_ack_1, ack => convolution3D_CP_1120_elements(6)); -- 
    rr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => type_cast_456_inst_req_0); -- 
    rr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(6), ack => RPIPE_maxpool_input_pipe_464_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Sample/ra
      -- 
    ra_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_0, ack => convolution3D_CP_1120_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_456_Update/ca
      -- 
    ca_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_1, ack => convolution3D_CP_1120_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_update_start_
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Update/cr
      -- 
    ra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_464_inst_ack_0, ack => convolution3D_CP_1120_elements(9)); -- 
    cr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(9), ack => RPIPE_maxpool_input_pipe_464_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_464_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Sample/rr
      -- 
    ca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_464_inst_ack_1, ack => convolution3D_CP_1120_elements(10)); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(10), ack => type_cast_468_inst_req_0); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(10), ack => RPIPE_maxpool_input_pipe_477_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Sample/ra
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_468_inst_ack_0, ack => convolution3D_CP_1120_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_468_Update/ca
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_468_inst_ack_1, ack => convolution3D_CP_1120_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_update_start_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Update/cr
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_477_inst_ack_0, ack => convolution3D_CP_1120_elements(13)); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(13), ack => RPIPE_maxpool_input_pipe_477_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_477_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Sample/rr
      -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_477_inst_ack_1, ack => convolution3D_CP_1120_elements(14)); -- 
    rr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => type_cast_481_inst_req_0); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => RPIPE_maxpool_input_pipe_489_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Sample/ra
      -- 
    ra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_0, ack => convolution3D_CP_1120_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_481_Update/ca
      -- 
    ca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_481_inst_ack_1, ack => convolution3D_CP_1120_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_update_start_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Update/cr
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_489_inst_ack_0, ack => convolution3D_CP_1120_elements(17)); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(17), ack => RPIPE_maxpool_input_pipe_489_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_489_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_sample_start_
      -- 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_489_inst_ack_1, ack => convolution3D_CP_1120_elements(18)); -- 
    rr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(18), ack => type_cast_493_inst_req_0); -- 
    rr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(18), ack => RPIPE_maxpool_input_pipe_502_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Sample/ra
      -- 
    ra_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_493_inst_ack_0, ack => convolution3D_CP_1120_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_493_Update/ca
      -- 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_493_inst_ack_1, ack => convolution3D_CP_1120_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_update_start_
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_sample_completed_
      -- 
    ra_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_502_inst_ack_0, ack => convolution3D_CP_1120_elements(21)); -- 
    cr_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(21), ack => RPIPE_maxpool_input_pipe_502_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_502_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Sample/$entry
      -- 
    ca_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_502_inst_ack_1, ack => convolution3D_CP_1120_elements(22)); -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => type_cast_506_inst_req_0); -- 
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => RPIPE_maxpool_input_pipe_514_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Sample/$exit
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_506_inst_ack_0, ack => convolution3D_CP_1120_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_506_Update/ca
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_506_inst_ack_1, ack => convolution3D_CP_1120_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_update_start_
      -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_514_inst_ack_0, ack => convolution3D_CP_1120_elements(25)); -- 
    cr_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(25), ack => RPIPE_maxpool_input_pipe_514_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_514_update_completed_
      -- 
    ca_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_514_inst_ack_1, ack => convolution3D_CP_1120_elements(26)); -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(26), ack => type_cast_518_inst_req_0); -- 
    rr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(26), ack => RPIPE_maxpool_input_pipe_527_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Sample/$exit
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_0, ack => convolution3D_CP_1120_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_518_Update/$exit
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_1, ack => convolution3D_CP_1120_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_update_start_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_sample_completed_
      -- 
    ra_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_527_inst_ack_0, ack => convolution3D_CP_1120_elements(29)); -- 
    cr_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(29), ack => RPIPE_maxpool_input_pipe_527_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_527_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Sample/rr
      -- 
    ca_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_527_inst_ack_1, ack => convolution3D_CP_1120_elements(30)); -- 
    rr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(30), ack => type_cast_531_inst_req_0); -- 
    rr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(30), ack => RPIPE_maxpool_input_pipe_539_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Sample/ra
      -- 
    ra_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_0, ack => convolution3D_CP_1120_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_531_update_completed_
      -- 
    ca_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_531_inst_ack_1, ack => convolution3D_CP_1120_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_update_start_
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Update/cr
      -- 
    ra_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_539_inst_ack_0, ack => convolution3D_CP_1120_elements(33)); -- 
    cr_1465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(33), ack => RPIPE_maxpool_input_pipe_539_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_539_Update/$exit
      -- 
    ca_1466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_539_inst_ack_1, ack => convolution3D_CP_1120_elements(34)); -- 
    rr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => type_cast_543_inst_req_0); -- 
    rr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(34), ack => RPIPE_maxpool_input_pipe_552_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_sample_completed_
      -- 
    ra_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_0, ack => convolution3D_CP_1120_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_543_update_completed_
      -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_1, ack => convolution3D_CP_1120_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_update_start_
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_sample_completed_
      -- 
    ra_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_552_inst_ack_0, ack => convolution3D_CP_1120_elements(37)); -- 
    cr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(37), ack => RPIPE_maxpool_input_pipe_552_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_552_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Sample/$entry
      -- 
    ca_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_552_inst_ack_1, ack => convolution3D_CP_1120_elements(38)); -- 
    rr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(38), ack => type_cast_556_inst_req_0); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(38), ack => RPIPE_maxpool_input_pipe_564_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Sample/ra
      -- 
    ra_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_0, ack => convolution3D_CP_1120_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_556_Update/ca
      -- 
    ca_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_1, ack => convolution3D_CP_1120_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_update_start_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Sample/$exit
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_564_inst_ack_0, ack => convolution3D_CP_1120_elements(41)); -- 
    cr_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(41), ack => RPIPE_maxpool_input_pipe_564_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_564_update_completed_
      -- 
    ca_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_564_inst_ack_1, ack => convolution3D_CP_1120_elements(42)); -- 
    rr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => type_cast_568_inst_req_0); -- 
    rr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => RPIPE_maxpool_input_pipe_577_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Sample/$exit
      -- 
    ra_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_568_inst_ack_0, ack => convolution3D_CP_1120_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_568_Update/$exit
      -- 
    ca_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_568_inst_ack_1, ack => convolution3D_CP_1120_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_update_start_
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Sample/$exit
      -- 
    ra_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_577_inst_ack_0, ack => convolution3D_CP_1120_elements(45)); -- 
    cr_1549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(45), ack => RPIPE_maxpool_input_pipe_577_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_577_update_completed_
      -- 
    ca_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_577_inst_ack_1, ack => convolution3D_CP_1120_elements(46)); -- 
    rr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(46), ack => type_cast_581_inst_req_0); -- 
    rr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(46), ack => RPIPE_maxpool_input_pipe_589_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Sample/ra
      -- 
    ra_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_581_inst_ack_0, ack => convolution3D_CP_1120_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_581_Update/$exit
      -- 
    ca_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_581_inst_ack_1, ack => convolution3D_CP_1120_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_update_start_
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_sample_completed_
      -- 
    ra_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_589_inst_ack_0, ack => convolution3D_CP_1120_elements(49)); -- 
    cr_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(49), ack => RPIPE_maxpool_input_pipe_589_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_589_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_sample_start_
      -- 
    ca_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_589_inst_ack_1, ack => convolution3D_CP_1120_elements(50)); -- 
    rr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => type_cast_593_inst_req_0); -- 
    rr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => RPIPE_maxpool_input_pipe_602_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Sample/ra
      -- 
    ra_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => convolution3D_CP_1120_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_593_Update/$exit
      -- 
    ca_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => convolution3D_CP_1120_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_update_start_
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Update/cr
      -- 
    ra_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_602_inst_ack_0, ack => convolution3D_CP_1120_elements(53)); -- 
    cr_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(53), ack => RPIPE_maxpool_input_pipe_602_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_602_Update/ca
      -- 
    ca_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_602_inst_ack_1, ack => convolution3D_CP_1120_elements(54)); -- 
    rr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(54), ack => type_cast_606_inst_req_0); -- 
    rr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(54), ack => RPIPE_maxpool_input_pipe_614_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Sample/ra
      -- 
    ra_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_0, ack => convolution3D_CP_1120_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_606_Update/ca
      -- 
    ca_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_1, ack => convolution3D_CP_1120_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_update_start_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Sample/ra
      -- 
    ra_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_614_inst_ack_0, ack => convolution3D_CP_1120_elements(57)); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(57), ack => RPIPE_maxpool_input_pipe_614_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_614_Update/$exit
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_614_inst_ack_1, ack => convolution3D_CP_1120_elements(58)); -- 
    rr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(58), ack => type_cast_618_inst_req_0); -- 
    rr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(58), ack => RPIPE_maxpool_input_pipe_627_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Sample/ra
      -- 
    ra_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_618_inst_ack_0, ack => convolution3D_CP_1120_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_618_Update/$exit
      -- 
    ca_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_618_inst_ack_1, ack => convolution3D_CP_1120_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_update_start_
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Update/cr
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Sample/$exit
      -- 
    ra_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_627_inst_ack_0, ack => convolution3D_CP_1120_elements(61)); -- 
    cr_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(61), ack => RPIPE_maxpool_input_pipe_627_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/RPIPE_maxpool_input_pipe_627_Update/$exit
      -- 
    ca_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_627_inst_ack_1, ack => convolution3D_CP_1120_elements(62)); -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(62), ack => type_cast_631_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_sample_completed_
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_0, ack => convolution3D_CP_1120_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_631_Update/ca
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_1, ack => convolution3D_CP_1120_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Sample/rr
      -- 
    rr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(65), ack => type_cast_640_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(12) & convolution3D_CP_1120_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Sample/ra
      -- 
    ra_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_640_inst_ack_0, ack => convolution3D_CP_1120_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_640_Update/$exit
      -- 
    ca_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_640_inst_ack_1, ack => convolution3D_CP_1120_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Sample/$entry
      -- 
    rr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(68), ack => type_cast_644_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(20) & convolution3D_CP_1120_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Sample/ra
      -- 
    ra_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_644_inst_ack_0, ack => convolution3D_CP_1120_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_644_Update/ca
      -- 
    ca_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_644_inst_ack_1, ack => convolution3D_CP_1120_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Sample/rr
      -- 
    rr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(71), ack => type_cast_660_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(4) & convolution3D_CP_1120_elements(8) & convolution3D_CP_1120_elements(67) & convolution3D_CP_1120_elements(70);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_sample_completed_
      -- 
    ra_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_0, ack => convolution3D_CP_1120_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/type_cast_660_Update/$exit
      -- 
    ca_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_1, ack => convolution3D_CP_1120_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/R_cmp321_669_place
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667__exit__
      -- CP-element group 74: 	 branch_block_stmt_436/if_stmt_668__entry__
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_440_to_assign_stmt_667/$exit
      -- 
    branch_req_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(74), ack => if_stmt_668_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(28) & convolution3D_CP_1120_elements(32) & convolution3D_CP_1120_elements(36) & convolution3D_CP_1120_elements(40) & convolution3D_CP_1120_elements(44) & convolution3D_CP_1120_elements(48) & convolution3D_CP_1120_elements(52) & convolution3D_CP_1120_elements(56) & convolution3D_CP_1120_elements(60) & convolution3D_CP_1120_elements(64) & convolution3D_CP_1120_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_436/entry_bbx_xnph323
      -- CP-element group 75: 	 branch_block_stmt_436/if_stmt_668_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/if_stmt_668_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_674__exit__
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743__entry__
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_update_start_
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_436/entry_bbx_xnph323_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/entry_bbx_xnph323_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_674_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_674_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_674_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/merge_stmt_674_PhiAck/dummy
      -- 
    if_choice_transition_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_668_branch_ack_1, ack => convolution3D_CP_1120_elements(75)); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_688_inst_req_0); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_688_inst_req_1); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_713_inst_req_0); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_704_inst_req_0); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_704_inst_req_1); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_713_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(75), ack => type_cast_723_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	274 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_436/if_stmt_668_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_436/if_stmt_668_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_940/$entry
      -- CP-element group 76: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/$entry
      -- 
    else_choice_transition_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_668_branch_ack_0, ack => convolution3D_CP_1120_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Sample/$exit
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_0, ack => convolution3D_CP_1120_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_688_Update/ca
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_1, ack => convolution3D_CP_1120_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Sample/$exit
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_0, ack => convolution3D_CP_1120_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_704_Update/ca
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_1, ack => convolution3D_CP_1120_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_sample_completed_
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_713_inst_ack_0, ack => convolution3D_CP_1120_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_713_Update/ca
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_713_inst_ack_1, ack => convolution3D_CP_1120_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Sample/rr
      -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(83), ack => type_cast_723_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(80) & convolution3D_CP_1120_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Sample/ra
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_723_inst_ack_0, ack => convolution3D_CP_1120_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/type_cast_723_Update/ca
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_723_inst_ack_1, ack => convolution3D_CP_1120_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	268 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743/$exit
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_679_to_assign_stmt_743__exit__
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_746/$entry
      -- CP-element group 86: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(78) & convolution3D_CP_1120_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	273 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Sample/ack
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_758_index_offset_ack_0, ack => convolution3D_CP_1120_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	273 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_request/req
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_758_index_offset_ack_1, ack => convolution3D_CP_1120_elements(88)); -- 
    req_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(88), ack => addr_of_759_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_request/ack
      -- 
    ack_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_759_final_reg_ack_0, ack => convolution3D_CP_1120_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	273 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_word_addrgen/root_register_ack
      -- 
    ack_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_759_final_reg_ack_1, ack => convolution3D_CP_1120_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	273 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_update_start_
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Update/cr
      -- 
    ra_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_762_inst_ack_0, ack => convolution3D_CP_1120_elements(91)); -- 
    cr_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(91), ack => RPIPE_maxpool_input_pipe_762_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Sample/rr
      -- 
    ca_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_762_inst_ack_1, ack => convolution3D_CP_1120_elements(92)); -- 
    rr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => type_cast_766_inst_req_0); -- 
    rr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => RPIPE_maxpool_input_pipe_775_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Sample/ra
      -- 
    ra_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_766_inst_ack_0, ack => convolution3D_CP_1120_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	273 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Update/ca
      -- 
    ca_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_766_inst_ack_1, ack => convolution3D_CP_1120_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_update_start_
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Update/cr
      -- 
    ra_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_775_inst_ack_0, ack => convolution3D_CP_1120_elements(95)); -- 
    cr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(95), ack => RPIPE_maxpool_input_pipe_775_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_775_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Sample/rr
      -- 
    ca_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_775_inst_ack_1, ack => convolution3D_CP_1120_elements(96)); -- 
    rr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(96), ack => type_cast_779_inst_req_0); -- 
    rr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(96), ack => RPIPE_maxpool_input_pipe_793_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Sample/ra
      -- 
    ra_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_0, ack => convolution3D_CP_1120_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	273 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Update/ca
      -- 
    ca_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_1, ack => convolution3D_CP_1120_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_update_start_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Update/cr
      -- 
    ra_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_793_inst_ack_0, ack => convolution3D_CP_1120_elements(99)); -- 
    cr_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(99), ack => RPIPE_maxpool_input_pipe_793_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_793_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Sample/rr
      -- 
    ca_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_793_inst_ack_1, ack => convolution3D_CP_1120_elements(100)); -- 
    rr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(100), ack => type_cast_797_inst_req_0); -- 
    rr_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(100), ack => RPIPE_maxpool_input_pipe_811_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Sample/ra
      -- 
    ra_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_0, ack => convolution3D_CP_1120_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	273 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Update/ca
      -- 
    ca_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_1, ack => convolution3D_CP_1120_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_update_start_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Update/cr
      -- 
    ra_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_811_inst_ack_0, ack => convolution3D_CP_1120_elements(103)); -- 
    cr_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(103), ack => RPIPE_maxpool_input_pipe_811_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_811_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Sample/rr
      -- 
    ca_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_811_inst_ack_1, ack => convolution3D_CP_1120_elements(104)); -- 
    rr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(104), ack => type_cast_815_inst_req_0); -- 
    rr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(104), ack => RPIPE_maxpool_input_pipe_829_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Sample/ra
      -- 
    ra_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_0, ack => convolution3D_CP_1120_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	273 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Update/ca
      -- 
    ca_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_1, ack => convolution3D_CP_1120_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_update_start_
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Update/cr
      -- 
    ra_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_829_inst_ack_0, ack => convolution3D_CP_1120_elements(107)); -- 
    cr_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(107), ack => RPIPE_maxpool_input_pipe_829_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_829_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Sample/rr
      -- 
    ca_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_829_inst_ack_1, ack => convolution3D_CP_1120_elements(108)); -- 
    rr_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(108), ack => type_cast_833_inst_req_0); -- 
    rr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(108), ack => RPIPE_maxpool_input_pipe_847_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Sample/ra
      -- 
    ra_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_0, ack => convolution3D_CP_1120_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	273 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Update/ca
      -- 
    ca_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_1, ack => convolution3D_CP_1120_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_update_start_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Update/cr
      -- 
    ra_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_847_inst_ack_0, ack => convolution3D_CP_1120_elements(111)); -- 
    cr_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(111), ack => RPIPE_maxpool_input_pipe_847_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_847_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Sample/rr
      -- 
    ca_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_847_inst_ack_1, ack => convolution3D_CP_1120_elements(112)); -- 
    rr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => type_cast_851_inst_req_0); -- 
    rr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => RPIPE_maxpool_input_pipe_865_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Sample/ra
      -- 
    ra_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => convolution3D_CP_1120_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	273 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Update/ca
      -- 
    ca_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => convolution3D_CP_1120_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_update_start_
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Update/cr
      -- 
    ra_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_865_inst_ack_0, ack => convolution3D_CP_1120_elements(115)); -- 
    cr_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(115), ack => RPIPE_maxpool_input_pipe_865_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_865_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Sample/rr
      -- 
    ca_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_865_inst_ack_1, ack => convolution3D_CP_1120_elements(116)); -- 
    rr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(116), ack => type_cast_869_inst_req_0); -- 
    rr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(116), ack => RPIPE_maxpool_input_pipe_883_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Sample/ra
      -- 
    ra_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_0, ack => convolution3D_CP_1120_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	273 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Update/ca
      -- 
    ca_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_1, ack => convolution3D_CP_1120_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_update_start_
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Update/cr
      -- 
    ra_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_883_inst_ack_0, ack => convolution3D_CP_1120_elements(119)); -- 
    cr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(119), ack => RPIPE_maxpool_input_pipe_883_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_883_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Sample/rr
      -- 
    ca_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_883_inst_ack_1, ack => convolution3D_CP_1120_elements(120)); -- 
    rr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(120), ack => type_cast_887_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Sample/ra
      -- 
    ra_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => convolution3D_CP_1120_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	273 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Update/ca
      -- 
    ca_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => convolution3D_CP_1120_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/ptr_deref_895_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/ptr_deref_895_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/ptr_deref_895_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/ptr_deref_895_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/word_access_start/word_0/rr
      -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(123), ack => ptr_deref_895_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(90) & convolution3D_CP_1120_elements(94) & convolution3D_CP_1120_elements(98) & convolution3D_CP_1120_elements(102) & convolution3D_CP_1120_elements(106) & convolution3D_CP_1120_elements(110) & convolution3D_CP_1120_elements(114) & convolution3D_CP_1120_elements(118) & convolution3D_CP_1120_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Sample/word_access_start/word_0/ra
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_895_store_0_ack_0, ack => convolution3D_CP_1120_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	273 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/word_access_complete/word_0/ca
      -- 
    ca_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_895_store_0_ack_1, ack => convolution3D_CP_1120_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	87 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908__exit__
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909__entry__
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_436/R_exitcond32_910_place
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_436/if_stmt_909_else_link/$entry
      -- 
    branch_req_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(126), ack => if_stmt_909_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(87) & convolution3D_CP_1120_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	275 
    -- CP-element group 127: 	276 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_915__exit__
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_922_to_assign_stmt_937__entry__
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_922_to_assign_stmt_937__exit__
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_915_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Update/cr
      -- CP-element group 127: 	 branch_block_stmt_436/if_stmt_909_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/if_stmt_909_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_922_to_assign_stmt_937/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_922_to_assign_stmt_937/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_915_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_915_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_436/merge_stmt_915_PhiReqMerge
      -- 
    if_choice_transition_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_909_branch_ack_1, ack => convolution3D_CP_1120_elements(127)); -- 
    rr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_943_inst_req_0); -- 
    cr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(127), ack => type_cast_943_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	269 
    -- CP-element group 128: 	270 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_436/if_stmt_909_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_436/if_stmt_909_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/$entry
      -- CP-element group 128: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/$entry
      -- 
    else_choice_transition_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_909_branch_ack_0, ack => convolution3D_CP_1120_elements(128)); -- 
    rr_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(128), ack => type_cast_752_inst_req_0); -- 
    cr_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(128), ack => type_cast_752_inst_req_1); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	279 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	298 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_436/if_stmt_960_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_436/if_stmt_960_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_436/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$entry
      -- 
    if_choice_transition_2157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_960_branch_ack_1, ack => convolution3D_CP_1120_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	279 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	280 
    -- CP-element group 130: 	281 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_966__exit__
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_972_to_assign_stmt_978__entry__
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_972_to_assign_stmt_978__exit__
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_966_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_966_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/if_stmt_960_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/if_stmt_960_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_972_to_assign_stmt_978/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_972_to_assign_stmt_978/$exit
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_966_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/merge_stmt_966_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/$entry
      -- 
    else_choice_transition_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_960_branch_ack_0, ack => convolution3D_CP_1120_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	293 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_update_start_
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Update/cr
      -- 
    ra_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1009_inst_ack_0, ack => convolution3D_CP_1120_elements(131)); -- 
    cr_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(131), ack => RPIPE_maxpool_input_pipe_1009_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Sample/rr
      -- 
    ca_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1009_inst_ack_1, ack => convolution3D_CP_1120_elements(132)); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(132), ack => type_cast_1013_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Sample/ra
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_0, ack => convolution3D_CP_1120_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	293 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Update/ca
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_1, ack => convolution3D_CP_1120_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	293 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Sample/ra
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1028_inst_ack_0, ack => convolution3D_CP_1120_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	293 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Update/ca
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1028_inst_ack_1, ack => convolution3D_CP_1120_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034__exit__
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035__entry__
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_436/R_cmpx_xi_1036_place
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/if_stmt_1035_else_link/$entry
      -- 
    branch_req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(137), ack => if_stmt_1035_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(134) & convolution3D_CP_1120_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	283 
    -- CP-element group 138: 	284 
    -- CP-element group 138: 	286 
    -- CP-element group 138: 	287 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_436/if_stmt_1035_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_436/if_stmt_1035_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- 
    if_choice_transition_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1035_branch_ack_1, ack => convolution3D_CP_1120_elements(138)); -- 
    rr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_994_inst_req_0); -- 
    cr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_994_inst_req_1); -- 
    cr_3448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_987_inst_req_1); -- 
    rr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => type_cast_987_inst_req_0); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	294 
    -- CP-element group 139: 	295 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/if_stmt_1035_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_436/if_stmt_1035_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1035_branch_ack_0, ack => convolution3D_CP_1120_elements(139)); -- 
    rr_3502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => type_cast_1045_inst_req_0); -- 
    cr_3507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => type_cast_1045_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	297 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Sample/ack
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1074_index_offset_ack_0, ack => convolution3D_CP_1120_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	297 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_request/req
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1074_index_offset_ack_1, ack => convolution3D_CP_1120_elements(141)); -- 
    req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(141), ack => addr_of_1075_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_request/ack
      -- 
    ack_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1075_final_reg_ack_0, ack => convolution3D_CP_1120_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	297 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/ptr_deref_1078_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/ptr_deref_1078_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/ptr_deref_1078_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/ptr_deref_1078_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/word_access_start/word_0/rr
      -- 
    ack_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1075_final_reg_ack_1, ack => convolution3D_CP_1120_elements(143)); -- 
    rr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(143), ack => ptr_deref_1078_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Sample/word_access_start/word_0/ra
      -- 
    ra_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1078_store_0_ack_0, ack => convolution3D_CP_1120_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	297 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/word_access_complete/word_0/ca
      -- 
    ca_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1078_store_0_ack_1, ack => convolution3D_CP_1120_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	298 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080__exit__
      -- CP-element group 146: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/$exit
      -- CP-element group 146: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- CP-element group 146: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(140) & convolution3D_CP_1120_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	298 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Sample/ra
      -- 
    ra_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_0, ack => convolution3D_CP_1120_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	298 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	155 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Update/ca
      -- 
    ca_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_1, ack => convolution3D_CP_1120_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	298 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Sample/ra
      -- 
    ra_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1089_inst_ack_0, ack => convolution3D_CP_1120_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	298 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Update/ca
      -- 
    ca_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1089_inst_ack_1, ack => convolution3D_CP_1120_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	298 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Sample/ra
      -- 
    ra_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1093_inst_ack_0, ack => convolution3D_CP_1120_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	298 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Update/ca
      -- 
    ca_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1093_inst_ack_1, ack => convolution3D_CP_1120_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	298 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Sample/ra
      -- 
    ra_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1097_inst_ack_0, ack => convolution3D_CP_1120_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	298 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Update/ca
      -- 
    ca_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1097_inst_ack_1, ack => convolution3D_CP_1120_elements(154)); -- 
    -- CP-element group 155:  branch  join  transition  place  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	148 
    -- CP-element group 155: 	150 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (10) 
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134__exit__
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135__entry__
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/$exit
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135_dead_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135_eval_test/$entry
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135_eval_test/$exit
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135_eval_test/branch_req
      -- CP-element group 155: 	 branch_block_stmt_436/R_cmp161317_1136_place
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135_if_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_436/if_stmt_1135_else_link/$entry
      -- 
    branch_req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(155), ack => if_stmt_1135_branch_req_0); -- 
    convolution3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(148) & convolution3D_CP_1120_elements(150) & convolution3D_CP_1120_elements(152) & convolution3D_CP_1120_elements(154);
      gj_convolution3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: 	159 
    -- CP-element group 156: 	160 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	162 
    -- CP-element group 156: 	163 
    -- CP-element group 156: 	164 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	168 
    -- CP-element group 156: 	170 
    -- CP-element group 156:  members (42) 
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1141__exit__
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212__entry__
      -- CP-element group 156: 	 branch_block_stmt_436/if_stmt_1135_if_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/if_stmt_1135_if_link/if_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_436/ifx_xend_bbx_xnph
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_update_start_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1141_PhiReqMerge
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1141_PhiAck/dummy
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1141_PhiAck/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/merge_stmt_1141_PhiAck/$entry
      -- CP-element group 156: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$entry
      -- 
    if_choice_transition_2401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1135_branch_ack_1, ack => convolution3D_CP_1120_elements(156)); -- 
    rr_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1156_inst_req_0); -- 
    cr_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1156_inst_req_1); -- 
    rr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1160_inst_req_0); -- 
    cr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1160_inst_req_1); -- 
    rr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1169_inst_req_0); -- 
    cr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1169_inst_req_1); -- 
    rr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1178_inst_req_0); -- 
    cr_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1178_inst_req_1); -- 
    cr_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1187_inst_req_1); -- 
    cr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(156), ack => type_cast_1192_inst_req_1); -- 
    -- CP-element group 157:  transition  place  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	308 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1409/$entry
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$entry
      -- CP-element group 157: 	 branch_block_stmt_436/if_stmt_1135_else_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_436/if_stmt_1135_else_link/else_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215
      -- CP-element group 157: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/$entry
      -- 
    else_choice_transition_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1135_branch_ack_0, ack => convolution3D_CP_1120_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Sample/ra
      -- 
    ra_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_0, ack => convolution3D_CP_1120_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	156 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	166 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1156_Update/ca
      -- 
    ca_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_1, ack => convolution3D_CP_1120_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	156 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Sample/ra
      -- 
    ra_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_0, ack => convolution3D_CP_1120_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	166 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1160_Update/ca
      -- 
    ca_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_1, ack => convolution3D_CP_1120_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	156 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Sample/ra
      -- 
    ra_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_0, ack => convolution3D_CP_1120_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	156 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1169_Update/ca
      -- 
    ca_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_1, ack => convolution3D_CP_1120_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Sample/ra
      -- 
    ra_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1178_inst_ack_0, ack => convolution3D_CP_1120_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1178_Update/ca
      -- 
    ca_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1178_inst_ack_1, ack => convolution3D_CP_1120_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	159 
    -- CP-element group 166: 	161 
    -- CP-element group 166: 	163 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Sample/rr
      -- 
    rr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(166), ack => type_cast_1187_inst_req_0); -- 
    convolution3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(159) & convolution3D_CP_1120_elements(161) & convolution3D_CP_1120_elements(163) & convolution3D_CP_1120_elements(165);
      gj_convolution3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Sample/ra
      -- 
    ra_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1187_inst_ack_0, ack => convolution3D_CP_1120_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	156 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1187_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Sample/rr
      -- 
    ca_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1187_inst_ack_1, ack => convolution3D_CP_1120_elements(168)); -- 
    rr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(168), ack => type_cast_1192_inst_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Sample/ra
      -- 
    ra_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_0, ack => convolution3D_CP_1120_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	156 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	299 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212__exit__
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/$exit
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_1147_to_assign_stmt_1212/type_cast_1192_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/$entry
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1215/$entry
      -- CP-element group 170: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- 
    ca_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_1, ack => convolution3D_CP_1120_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	304 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_sample_complete
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1227_index_offset_ack_0, ack => convolution3D_CP_1120_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	304 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_request/req
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_offset_calculated
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Update/$exit
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1227_index_offset_ack_1, ack => convolution3D_CP_1120_elements(172)); -- 
    req_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(172), ack => addr_of_1228_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_request/ack
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_sample_completed_
      -- 
    ack_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1228_final_reg_ack_0, ack => convolution3D_CP_1120_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	304 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_complete/ack
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_word_addrgen/root_register_ack
      -- 
    ack_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1228_final_reg_ack_1, ack => convolution3D_CP_1120_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	304 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_update_start_
      -- 
    ra_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1231_inst_ack_0, ack => convolution3D_CP_1120_elements(175)); -- 
    cr_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(175), ack => RPIPE_maxpool_input_pipe_1231_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Sample/$entry
      -- 
    ca_2557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1231_inst_ack_1, ack => convolution3D_CP_1120_elements(176)); -- 
    rr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(176), ack => type_cast_1235_inst_req_0); -- 
    rr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(176), ack => RPIPE_maxpool_input_pipe_1244_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Sample/$exit
      -- 
    ra_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_0, ack => convolution3D_CP_1120_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	304 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_update_completed_
      -- 
    ca_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_1, ack => convolution3D_CP_1120_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_update_start_
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_sample_completed_
      -- 
    ra_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1244_inst_ack_0, ack => convolution3D_CP_1120_elements(179)); -- 
    cr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(179), ack => RPIPE_maxpool_input_pipe_1244_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1244_update_completed_
      -- 
    ca_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1244_inst_ack_1, ack => convolution3D_CP_1120_elements(180)); -- 
    rr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => type_cast_1248_inst_req_0); -- 
    rr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => RPIPE_maxpool_input_pipe_1262_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_sample_completed_
      -- 
    ra_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_0, ack => convolution3D_CP_1120_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	304 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_update_completed_
      -- 
    ca_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_1, ack => convolution3D_CP_1120_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_update_start_
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Update/$entry
      -- 
    ra_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1262_inst_ack_0, ack => convolution3D_CP_1120_elements(183)); -- 
    cr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(183), ack => RPIPE_maxpool_input_pipe_1262_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1262_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Sample/$entry
      -- 
    ca_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1262_inst_ack_1, ack => convolution3D_CP_1120_elements(184)); -- 
    rr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(184), ack => type_cast_1266_inst_req_0); -- 
    rr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(184), ack => RPIPE_maxpool_input_pipe_1280_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Sample/$exit
      -- 
    ra_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_0, ack => convolution3D_CP_1120_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	304 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_update_completed_
      -- 
    ca_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_1, ack => convolution3D_CP_1120_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_update_start_
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_sample_completed_
      -- 
    ra_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1280_inst_ack_0, ack => convolution3D_CP_1120_elements(187)); -- 
    cr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => RPIPE_maxpool_input_pipe_1280_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1280_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_sample_start_
      -- 
    ca_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1280_inst_ack_1, ack => convolution3D_CP_1120_elements(188)); -- 
    rr_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(188), ack => type_cast_1284_inst_req_0); -- 
    rr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(188), ack => RPIPE_maxpool_input_pipe_1298_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Sample/ra
      -- 
    ra_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_0, ack => convolution3D_CP_1120_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	304 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Update/$exit
      -- 
    ca_2655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_1, ack => convolution3D_CP_1120_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_update_start_
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_sample_completed_
      -- 
    ra_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1298_inst_ack_0, ack => convolution3D_CP_1120_elements(191)); -- 
    cr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(191), ack => RPIPE_maxpool_input_pipe_1298_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1298_Update/ca
      -- 
    ca_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1298_inst_ack_1, ack => convolution3D_CP_1120_elements(192)); -- 
    rr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(192), ack => type_cast_1302_inst_req_0); -- 
    rr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(192), ack => RPIPE_maxpool_input_pipe_1316_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_sample_completed_
      -- 
    ra_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_0, ack => convolution3D_CP_1120_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	304 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_update_completed_
      -- 
    ca_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_1, ack => convolution3D_CP_1120_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_update_start_
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Update/cr
      -- 
    ra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1316_inst_ack_0, ack => convolution3D_CP_1120_elements(195)); -- 
    cr_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(195), ack => RPIPE_maxpool_input_pipe_1316_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1316_Update/$exit
      -- 
    ca_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1316_inst_ack_1, ack => convolution3D_CP_1120_elements(196)); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(196), ack => type_cast_1320_inst_req_0); -- 
    rr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(196), ack => RPIPE_maxpool_input_pipe_1334_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_sample_completed_
      -- 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => convolution3D_CP_1120_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	304 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_update_completed_
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => convolution3D_CP_1120_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Update/cr
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_update_start_
      -- 
    ra_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1334_inst_ack_0, ack => convolution3D_CP_1120_elements(199)); -- 
    cr_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(199), ack => RPIPE_maxpool_input_pipe_1334_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1334_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Sample/rr
      -- 
    ca_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1334_inst_ack_1, ack => convolution3D_CP_1120_elements(200)); -- 
    rr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(200), ack => type_cast_1338_inst_req_0); -- 
    rr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(200), ack => RPIPE_maxpool_input_pipe_1352_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Sample/$exit
      -- 
    ra_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_0, ack => convolution3D_CP_1120_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	304 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Update/ca
      -- 
    ca_2739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_1, ack => convolution3D_CP_1120_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_update_start_
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Update/cr
      -- 
    ra_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1352_inst_ack_0, ack => convolution3D_CP_1120_elements(203)); -- 
    cr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(203), ack => RPIPE_maxpool_input_pipe_1352_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1352_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Sample/rr
      -- 
    ca_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1352_inst_ack_1, ack => convolution3D_CP_1120_elements(204)); -- 
    rr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(204), ack => type_cast_1356_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Sample/ra
      -- 
    ra_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_0, ack => convolution3D_CP_1120_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	304 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Update/ca
      -- 
    ca_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_1, ack => convolution3D_CP_1120_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/ptr_deref_1364_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/ptr_deref_1364_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/ptr_deref_1364_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/ptr_deref_1364_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/word_access_start/word_0/rr
      -- 
    rr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(207), ack => ptr_deref_1364_store_0_req_0); -- 
    convolution3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(174) & convolution3D_CP_1120_elements(178) & convolution3D_CP_1120_elements(182) & convolution3D_CP_1120_elements(186) & convolution3D_CP_1120_elements(190) & convolution3D_CP_1120_elements(194) & convolution3D_CP_1120_elements(198) & convolution3D_CP_1120_elements(202) & convolution3D_CP_1120_elements(206);
      gj_convolution3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Sample/word_access_start/word_0/ra
      -- 
    ra_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1364_store_0_ack_0, ack => convolution3D_CP_1120_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	304 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/word_access_complete/word_0/ca
      -- 
    ca_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1364_store_0_ack_1, ack => convolution3D_CP_1120_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	171 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_436/R_exitcond_1379_place
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377__exit__
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378__entry__
      -- CP-element group 210: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/$exit
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1378_else_link/$entry
      -- 
    branch_req_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => if_stmt_1378_branch_req_0); -- 
    convolution3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(171) & convolution3D_CP_1120_elements(209);
      gj_convolution3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	305 
    -- CP-element group 211: 	306 
    -- CP-element group 211:  members (24) 
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1384_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1384__exit__
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1391_to_assign_stmt_1406__entry__
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1391_to_assign_stmt_1406__exit__
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 211: 	 branch_block_stmt_436/if_stmt_1378_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/if_stmt_1378_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1391_to_assign_stmt_1406/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/assign_stmt_1391_to_assign_stmt_1406/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Update/cr
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1384_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1384_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/merge_stmt_1384_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- 
    if_choice_transition_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1378_branch_ack_1, ack => convolution3D_CP_1120_elements(211)); -- 
    cr_3615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => type_cast_1412_inst_req_1); -- 
    rr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => type_cast_1412_inst_req_0); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	300 
    -- CP-element group 212: 	301 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Update/cr
      -- CP-element group 212: 	 branch_block_stmt_436/if_stmt_1378_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_436/if_stmt_1378_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/$entry
      -- CP-element group 212: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- 
    else_choice_transition_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1378_branch_ack_0, ack => convolution3D_CP_1120_elements(212)); -- 
    rr_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_1221_inst_req_0); -- 
    cr_3572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(212), ack => type_cast_1221_inst_req_1); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	310 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	329 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_436/if_stmt_1429_if_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_436/if_stmt_1429_if_link/if_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_436/forx_xend215_ifx_xend227
      -- CP-element group 213: 	 branch_block_stmt_436/forx_xend215_ifx_xend227_PhiReq/$exit
      -- CP-element group 213: 	 branch_block_stmt_436/forx_xend215_ifx_xend227_PhiReq/$entry
      -- 
    if_choice_transition_2855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1429_branch_ack_1, ack => convolution3D_CP_1120_elements(213)); -- 
    -- CP-element group 214:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	310 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (18) 
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1435__exit__
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451__entry__
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1435_PhiReqMerge
      -- CP-element group 214: 	 branch_block_stmt_436/forx_xend215_bbx_xnphx_xi294_PhiReq/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/forx_xend215_bbx_xnphx_xi294_PhiReq/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1435_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1435_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1429_else_link/$exit
      -- CP-element group 214: 	 branch_block_stmt_436/if_stmt_1429_else_link/else_choice_transition
      -- CP-element group 214: 	 branch_block_stmt_436/forx_xend215_bbx_xnphx_xi294
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_update_start_
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Update/cr
      -- CP-element group 214: 	 branch_block_stmt_436/merge_stmt_1435_PhiAck/dummy
      -- 
    else_choice_transition_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1429_branch_ack_0, ack => convolution3D_CP_1120_elements(214)); -- 
    rr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(214), ack => type_cast_1444_inst_req_0); -- 
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(214), ack => type_cast_1444_inst_req_1); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Sample/ra
      -- 
    ra_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1444_inst_ack_0, ack => convolution3D_CP_1120_elements(215)); -- 
    -- CP-element group 216:  fork  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	311 
    -- CP-element group 216: 	312 
    -- CP-element group 216:  members (11) 
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451__exit__
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1441_to_assign_stmt_1451/type_cast_1444_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/$entry
      -- CP-element group 216: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/$entry
      -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1444_inst_ack_1, ack => convolution3D_CP_1120_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	324 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_update_start_
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Update/cr
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1482_inst_ack_0, ack => convolution3D_CP_1120_elements(217)); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(217), ack => RPIPE_maxpool_input_pipe_1482_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Sample/rr
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1482_inst_ack_1, ack => convolution3D_CP_1120_elements(218)); -- 
    rr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(218), ack => type_cast_1486_inst_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Sample/ra
      -- 
    ra_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1486_inst_ack_0, ack => convolution3D_CP_1120_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	324 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Update/ca
      -- 
    ca_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1486_inst_ack_1, ack => convolution3D_CP_1120_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	324 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Sample/ra
      -- 
    ra_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1501_inst_ack_0, ack => convolution3D_CP_1120_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	324 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Update/ca
      -- 
    ca_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1501_inst_ack_1, ack => convolution3D_CP_1120_elements(222)); -- 
    -- CP-element group 223:  branch  join  transition  place  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507__exit__
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508__entry__
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/$exit
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508_dead_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508_eval_test/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508_eval_test/$exit
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508_eval_test/branch_req
      -- CP-element group 223: 	 branch_block_stmt_436/R_cmpx_xi302_1509_place
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508_if_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_436/if_stmt_1508_else_link/$entry
      -- 
    branch_req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(223), ack => if_stmt_1508_branch_req_0); -- 
    convolution3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(220) & convolution3D_CP_1120_elements(222);
      gj_convolution3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	314 
    -- CP-element group 224: 	315 
    -- CP-element group 224: 	317 
    -- CP-element group 224: 	318 
    -- CP-element group 224:  members (20) 
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/if_stmt_1508_if_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_436/if_stmt_1508_if_link/if_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Update/$entry
      -- 
    if_choice_transition_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1508_branch_ack_1, ack => convolution3D_CP_1120_elements(224)); -- 
    rr_3683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1460_inst_req_0); -- 
    cr_3711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1467_inst_req_1); -- 
    rr_3706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1467_inst_req_0); -- 
    cr_3688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(224), ack => type_cast_1460_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	325 
    -- CP-element group 225: 	326 
    -- CP-element group 225:  members (12) 
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Update/cr
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/if_stmt_1508_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_436/if_stmt_1508_else_link/else_choice_transition
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 225: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/$entry
      -- 
    else_choice_transition_2940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1508_branch_ack_0, ack => convolution3D_CP_1120_elements(225)); -- 
    cr_3747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(225), ack => type_cast_1518_inst_req_1); -- 
    rr_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(225), ack => type_cast_1518_inst_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	328 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	232 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_sample_complete
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Sample/ack
      -- 
    ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1547_index_offset_ack_0, ack => convolution3D_CP_1120_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	328 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (11) 
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_offset_calculated
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Update/ack
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_base_plus_offset/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_base_plus_offset/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_base_plus_offset/sum_rename_req
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_base_plus_offset/sum_rename_ack
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_request/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_request/req
      -- 
    ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1547_index_offset_ack_1, ack => convolution3D_CP_1120_elements(227)); -- 
    req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(227), ack => addr_of_1548_final_reg_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_request/$exit
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_request/ack
      -- 
    ack_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1548_final_reg_ack_0, ack => convolution3D_CP_1120_elements(228)); -- 
    -- CP-element group 229:  join  fork  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	328 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (28) 
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_complete/ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_word_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_address_resized
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_addr_resize/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_addr_resize/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_addr_resize/base_resize_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_addr_resize/base_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_word_addrgen/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_word_addrgen/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_word_addrgen/root_register_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_word_addrgen/root_register_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/ptr_deref_1551_Split/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/ptr_deref_1551_Split/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/ptr_deref_1551_Split/split_req
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/ptr_deref_1551_Split/split_ack
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/word_access_start/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/word_access_start/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/word_access_start/word_0/rr
      -- 
    ack_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1548_final_reg_ack_1, ack => convolution3D_CP_1120_elements(229)); -- 
    rr_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(229), ack => ptr_deref_1551_store_0_req_0); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Sample/word_access_start/word_0/ra
      -- 
    ra_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1551_store_0_ack_0, ack => convolution3D_CP_1120_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	328 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/word_access_complete/word_0/ca
      -- 
    ca_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1551_store_0_ack_1, ack => convolution3D_CP_1120_elements(231)); -- 
    -- CP-element group 232:  join  transition  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	226 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	329 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553__exit__
      -- CP-element group 232: 	 branch_block_stmt_436/getRemainingElementsx_xexit311_ifx_xend227
      -- CP-element group 232: 	 branch_block_stmt_436/getRemainingElementsx_xexit311_ifx_xend227_PhiReq/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/getRemainingElementsx_xexit311_ifx_xend227_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(226) & convolution3D_CP_1120_elements(231);
      gj_convolution3D_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	329 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Sample/cra
      -- 
    cra_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1558_call_ack_0, ack => convolution3D_CP_1120_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	329 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	237 
    -- CP-element group 234: 	241 
    -- CP-element group 234: 	242 
    -- CP-element group 234: 	243 
    -- CP-element group 234: 	244 
    -- CP-element group 234: 	245 
    -- CP-element group 234: 	246 
    -- CP-element group 234:  members (31) 
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1558__exit__
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626__entry__
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1558/$exit
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Update/cca
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_update_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_update_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_update_start_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Update/cr
      -- 
    cca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1558_call_ack_1, ack => convolution3D_CP_1120_elements(234)); -- 
    req_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => WPIPE_num_out_pipe_1570_inst_req_0); -- 
    req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => WPIPE_maxpool_output_pipe_1573_inst_req_0); -- 
    rr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1601_inst_req_0); -- 
    cr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1601_inst_req_1); -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1611_inst_req_0); -- 
    cr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1611_inst_req_1); -- 
    rr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1620_inst_req_0); -- 
    cr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(234), ack => type_cast_1620_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_update_start_
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Update/req
      -- 
    ack_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1570_inst_ack_0, ack => convolution3D_CP_1120_elements(235)); -- 
    req_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(235), ack => WPIPE_num_out_pipe_1570_inst_req_1); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	247 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_num_out_pipe_1570_Update/ack
      -- 
    ack_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1570_inst_ack_1, ack => convolution3D_CP_1120_elements(236)); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	234 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_update_start_
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Update/req
      -- 
    ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1573_inst_ack_0, ack => convolution3D_CP_1120_elements(237)); -- 
    req_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(237), ack => WPIPE_maxpool_output_pipe_1573_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1573_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Sample/req
      -- 
    ack_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1573_inst_ack_1, ack => convolution3D_CP_1120_elements(238)); -- 
    req_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(238), ack => WPIPE_maxpool_output_pipe_1577_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_update_start_
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Update/req
      -- 
    ack_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1577_inst_ack_0, ack => convolution3D_CP_1120_elements(239)); -- 
    req_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(239), ack => WPIPE_maxpool_output_pipe_1577_inst_req_1); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	247 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/WPIPE_maxpool_output_pipe_1577_Update/ack
      -- 
    ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1577_inst_ack_1, ack => convolution3D_CP_1120_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	234 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Sample/ra
      -- 
    ra_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_0, ack => convolution3D_CP_1120_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	234 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	247 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1601_Update/ca
      -- 
    ca_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_1, ack => convolution3D_CP_1120_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	234 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Sample/ra
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_0, ack => convolution3D_CP_1120_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	234 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	247 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1611_Update/ca
      -- 
    ca_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_1, ack => convolution3D_CP_1120_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	234 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Sample/ra
      -- 
    ra_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1620_inst_ack_0, ack => convolution3D_CP_1120_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	234 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/type_cast_1620_Update/ca
      -- 
    ca_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1620_inst_ack_1, ack => convolution3D_CP_1120_elements(246)); -- 
    -- CP-element group 247:  join  transition  place  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	236 
    -- CP-element group 247: 	240 
    -- CP-element group 247: 	242 
    -- CP-element group 247: 	244 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	330 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626__exit__
      -- CP-element group 247: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody
      -- CP-element group 247: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1629/$entry
      -- CP-element group 247: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1564_to_assign_stmt_1626/$exit
      -- CP-element group 247: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/$entry
      -- 
    convolution3D_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(236) & convolution3D_CP_1120_elements(240) & convolution3D_CP_1120_elements(242) & convolution3D_CP_1120_elements(244) & convolution3D_CP_1120_elements(246);
      gj_convolution3D_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	335 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Sample/ra
      -- 
    ra_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1649_inst_ack_0, ack => convolution3D_CP_1120_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	335 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Update/ca
      -- 
    ca_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1649_inst_ack_1, ack => convolution3D_CP_1120_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	335 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Sample/ra
      -- 
    ra_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1653_inst_ack_0, ack => convolution3D_CP_1120_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	335 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Update/ca
      -- 
    ca_3176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1653_inst_ack_1, ack => convolution3D_CP_1120_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Sample/crr
      -- 
    crr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(252), ack => call_stmt_1657_call_req_0); -- 
    convolution3D_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(249) & convolution3D_CP_1120_elements(251);
      gj_convolution3D_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Sample/cra
      -- 
    cra_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1657_call_ack_0, ack => convolution3D_CP_1120_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	335 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	257 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Update/cca
      -- 
    cca_3190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1657_call_ack_1, ack => convolution3D_CP_1120_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	335 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Sample/cra
      -- 
    cra_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1664_call_ack_0, ack => convolution3D_CP_1120_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	335 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Update/cca
      -- 
    cca_3204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1664_call_ack_1, ack => convolution3D_CP_1120_elements(256)); -- 
    -- CP-element group 257:  branch  join  transition  place  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	254 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (10) 
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675__exit__
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676__entry__
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/$exit
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676_dead_link/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676_eval_test/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676_eval_test/$exit
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676_eval_test/branch_req
      -- CP-element group 257: 	 branch_block_stmt_436/R_exitcond5_1677_place
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676_if_link/$entry
      -- CP-element group 257: 	 branch_block_stmt_436/if_stmt_1676_else_link/$entry
      -- 
    branch_req_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(257), ack => if_stmt_1676_branch_req_0); -- 
    convolution3D_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(254) & convolution3D_CP_1120_elements(256);
      gj_convolution3D_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	261 
    -- CP-element group 258:  members (18) 
      -- CP-element group 258: 	 branch_block_stmt_436/merge_stmt_1682__exit__
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687__entry__
      -- CP-element group 258: 	 branch_block_stmt_436/merge_stmt_1682_PhiReqMerge
      -- CP-element group 258: 	 branch_block_stmt_436/if_stmt_1676_if_link/$exit
      -- CP-element group 258: 	 branch_block_stmt_436/if_stmt_1676_if_link/if_choice_transition
      -- CP-element group 258: 	 branch_block_stmt_436/whilex_xbody_whilex_xend
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/$entry
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_update_start_
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Sample/rr
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Update/cr
      -- CP-element group 258: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 258: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 258: 	 branch_block_stmt_436/merge_stmt_1682_PhiAck/$entry
      -- CP-element group 258: 	 branch_block_stmt_436/merge_stmt_1682_PhiAck/$exit
      -- CP-element group 258: 	 branch_block_stmt_436/merge_stmt_1682_PhiAck/dummy
      -- 
    if_choice_transition_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1676_branch_ack_1, ack => convolution3D_CP_1120_elements(258)); -- 
    rr_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(258), ack => type_cast_1686_inst_req_0); -- 
    cr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(258), ack => type_cast_1686_inst_req_1); -- 
    -- CP-element group 259:  fork  transition  place  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	331 
    -- CP-element group 259: 	332 
    -- CP-element group 259:  members (12) 
      -- CP-element group 259: 	 branch_block_stmt_436/if_stmt_1676_else_link/$exit
      -- CP-element group 259: 	 branch_block_stmt_436/if_stmt_1676_else_link/else_choice_transition
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1676_branch_ack_0, ack => convolution3D_CP_1120_elements(259)); -- 
    rr_3795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => type_cast_1632_inst_req_0); -- 
    cr_3800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(259), ack => type_cast_1632_inst_req_1); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Sample/ra
      -- 
    ra_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_0, ack => convolution3D_CP_1120_elements(260)); -- 
    -- CP-element group 261:  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	258 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	265 
    -- CP-element group 261:  members (16) 
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1687__exit__
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703__entry__
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1687/$exit
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1687/type_cast_1686_Update/ca
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_update_start_
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Sample/crr
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Update/ccr
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_update_start_
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Update/cr
      -- 
    ca_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_1, ack => convolution3D_CP_1120_elements(261)); -- 
    crr_3251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => call_stmt_1690_call_req_0); -- 
    ccr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => call_stmt_1690_call_req_1); -- 
    cr_3270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => type_cast_1694_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Sample/cra
      -- 
    cra_3252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1690_call_ack_0, ack => convolution3D_CP_1120_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/call_stmt_1690_Update/cca
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Sample/rr
      -- 
    cca_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1690_call_ack_1, ack => convolution3D_CP_1120_elements(263)); -- 
    rr_3265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(263), ack => type_cast_1694_inst_req_0); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Sample/ra
      -- 
    ra_3266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_0, ack => convolution3D_CP_1120_elements(264)); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	261 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/type_cast_1694_Update/ca
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Sample/req
      -- 
    ca_3271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_1, ack => convolution3D_CP_1120_elements(265)); -- 
    req_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(265), ack => WPIPE_elapsed_time_pipe_1701_inst_req_0); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_update_start_
      -- CP-element group 266: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Sample/ack
      -- CP-element group 266: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Update/req
      -- 
    ack_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1701_inst_ack_0, ack => convolution3D_CP_1120_elements(266)); -- 
    req_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(266), ack => WPIPE_elapsed_time_pipe_1701_inst_req_1); -- 
    -- CP-element group 267:  transition  place  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (16) 
      -- CP-element group 267: 	 $exit
      -- CP-element group 267: 	 branch_block_stmt_436/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/branch_block_stmt_436__exit__
      -- CP-element group 267: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703__exit__
      -- CP-element group 267: 	 branch_block_stmt_436/return__
      -- CP-element group 267: 	 branch_block_stmt_436/merge_stmt_1706__exit__
      -- CP-element group 267: 	 branch_block_stmt_436/merge_stmt_1706_PhiReqMerge
      -- CP-element group 267: 	 branch_block_stmt_436/merge_stmt_1706_PhiAck/$entry
      -- CP-element group 267: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/call_stmt_1690_to_assign_stmt_1703/WPIPE_elapsed_time_pipe_1701_Update/ack
      -- CP-element group 267: 	 branch_block_stmt_436/return___PhiReq/$entry
      -- CP-element group 267: 	 branch_block_stmt_436/return___PhiReq/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/merge_stmt_1706_PhiAck/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/merge_stmt_1706_PhiAck/dummy
      -- 
    ack_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1701_inst_ack_1, ack => convolution3D_CP_1120_elements(267)); -- 
    -- CP-element group 268:  transition  output  delay-element  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	86 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	272 
    -- CP-element group 268:  members (5) 
      -- CP-element group 268: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/$exit
      -- CP-element group 268: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_746/$exit
      -- CP-element group 268: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/$exit
      -- CP-element group 268: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_750_konst_delay_trans
      -- CP-element group 268: 	 branch_block_stmt_436/bbx_xnph323_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_req
      -- 
    phi_stmt_746_req_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_746_req_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(268), ack => phi_stmt_746_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(268) is a control-delay.
    cp_element_268_delay: control_delay_element  generic map(name => " 268_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(86), ack => convolution3D_CP_1120_elements(268), clk => clk, reset =>reset);
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	128 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (2) 
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Sample/ra
      -- 
    ra_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_0, ack => convolution3D_CP_1120_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	128 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/Update/ca
      -- 
    ca_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_1, ack => convolution3D_CP_1120_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_req
      -- CP-element group 271: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_746/phi_stmt_746_sources/type_cast_752/SplitProtocol/$exit
      -- 
    phi_stmt_746_req_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_746_req_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(271), ack => phi_stmt_746_req_1); -- 
    convolution3D_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(269) & convolution3D_CP_1120_elements(270);
      gj_convolution3D_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  merge  transition  place  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	268 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (2) 
      -- CP-element group 272: 	 branch_block_stmt_436/merge_stmt_745_PhiAck/$entry
      -- CP-element group 272: 	 branch_block_stmt_436/merge_stmt_745_PhiReqMerge
      -- 
    convolution3D_CP_1120_elements(272) <= OrReduce(convolution3D_CP_1120_elements(268) & convolution3D_CP_1120_elements(271));
    -- CP-element group 273:  fork  transition  place  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	87 
    -- CP-element group 273: 	88 
    -- CP-element group 273: 	90 
    -- CP-element group 273: 	91 
    -- CP-element group 273: 	94 
    -- CP-element group 273: 	98 
    -- CP-element group 273: 	102 
    -- CP-element group 273: 	106 
    -- CP-element group 273: 	110 
    -- CP-element group 273: 	114 
    -- CP-element group 273: 	118 
    -- CP-element group 273: 	122 
    -- CP-element group 273: 	125 
    -- CP-element group 273:  members (56) 
      -- CP-element group 273: 	 branch_block_stmt_436/merge_stmt_745__exit__
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908__entry__
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_resized_1
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_scaled_1
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_computed_1
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_resize_1/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_resize_1/$exit
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_resize_1/index_resize_req
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_resize_1/index_resize_ack
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_scale_1/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_scale_1/$exit
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_scale_1/scale_rename_req
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_index_scale_1/scale_rename_ack
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_update_start
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Sample/req
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/array_obj_ref_758_final_index_sum_regn_Update/req
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_complete/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/addr_of_759_complete/req
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_sample_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/RPIPE_maxpool_input_pipe_762_Sample/rr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_766_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_779_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_797_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_815_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_833_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_851_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_869_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/type_cast_887_Update/cr
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_update_start_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/word_access_complete/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/word_access_complete/word_0/$entry
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_760_to_assign_stmt_908/ptr_deref_895_Update/word_access_complete/word_0/cr
      -- CP-element group 273: 	 branch_block_stmt_436/merge_stmt_745_PhiAck/$exit
      -- CP-element group 273: 	 branch_block_stmt_436/merge_stmt_745_PhiAck/phi_stmt_746_ack
      -- 
    phi_stmt_746_ack_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_746_ack_0, ack => convolution3D_CP_1120_elements(273)); -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => array_obj_ref_758_index_offset_req_0); -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => array_obj_ref_758_index_offset_req_1); -- 
    req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => addr_of_759_final_reg_req_1); -- 
    rr_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => RPIPE_maxpool_input_pipe_762_inst_req_0); -- 
    cr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_766_inst_req_1); -- 
    cr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_779_inst_req_1); -- 
    cr_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_797_inst_req_1); -- 
    cr_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_815_inst_req_1); -- 
    cr_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_833_inst_req_1); -- 
    cr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_851_inst_req_1); -- 
    cr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_869_inst_req_1); -- 
    cr_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => type_cast_887_inst_req_1); -- 
    cr_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(273), ack => ptr_deref_895_store_0_req_1); -- 
    -- CP-element group 274:  transition  output  delay-element  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	76 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	278 
    -- CP-element group 274:  members (5) 
      -- CP-element group 274: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$exit
      -- CP-element group 274: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_940/$exit
      -- CP-element group 274: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_req
      -- CP-element group 274: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_946_konst_delay_trans
      -- CP-element group 274: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/$exit
      -- 
    phi_stmt_940_req_3362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_940_req_3362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(274), ack => phi_stmt_940_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(274) is a control-delay.
    cp_element_274_delay: control_delay_element  generic map(name => " 274_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(76), ack => convolution3D_CP_1120_elements(274), clk => clk, reset =>reset);
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	127 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (2) 
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Sample/ra
      -- 
    ra_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_943_inst_ack_0, ack => convolution3D_CP_1120_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	127 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (2) 
      -- CP-element group 276: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/Update/ca
      -- 
    ca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_943_inst_ack_1, ack => convolution3D_CP_1120_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/type_cast_943/SplitProtocol/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_req
      -- CP-element group 277: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/phi_stmt_940_sources/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_940/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_940_req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_940_req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(277), ack => phi_stmt_940_req_0); -- 
    convolution3D_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(275) & convolution3D_CP_1120_elements(276);
      gj_convolution3D_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  merge  transition  place  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	274 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_436/merge_stmt_939_PhiAck/$entry
      -- CP-element group 278: 	 branch_block_stmt_436/merge_stmt_939_PhiReqMerge
      -- 
    convolution3D_CP_1120_elements(278) <= OrReduce(convolution3D_CP_1120_elements(274) & convolution3D_CP_1120_elements(277));
    -- CP-element group 279:  branch  transition  place  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	129 
    -- CP-element group 279: 	130 
    -- CP-element group 279:  members (15) 
      -- CP-element group 279: 	 branch_block_stmt_436/merge_stmt_939__exit__
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_953_to_assign_stmt_959__entry__
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_953_to_assign_stmt_959__exit__
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960__entry__
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_953_to_assign_stmt_959/$entry
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_953_to_assign_stmt_959/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960_dead_link/$entry
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960_eval_test/$entry
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960_eval_test/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960_eval_test/branch_req
      -- CP-element group 279: 	 branch_block_stmt_436/R_tobool_961_place
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960_if_link/$entry
      -- CP-element group 279: 	 branch_block_stmt_436/if_stmt_960_else_link/$entry
      -- CP-element group 279: 	 branch_block_stmt_436/merge_stmt_939_PhiAck/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/merge_stmt_939_PhiAck/phi_stmt_940_ack
      -- 
    phi_stmt_940_ack_3393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_940_ack_0, ack => convolution3D_CP_1120_elements(279)); -- 
    branch_req_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(279), ack => if_stmt_960_branch_req_0); -- 
    -- CP-element group 280:  transition  output  delay-element  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	130 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (4) 
      -- CP-element group 280: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_req
      -- CP-element group 280: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_985_konst_delay_trans
      -- CP-element group 280: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/$exit
      -- CP-element group 280: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/$exit
      -- 
    phi_stmt_981_req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_981_req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(280), ack => phi_stmt_981_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(280) is a control-delay.
    cp_element_280_delay: control_delay_element  generic map(name => " 280_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(130), ack => convolution3D_CP_1120_elements(280), clk => clk, reset =>reset);
    -- CP-element group 281:  transition  output  delay-element  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	130 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (4) 
      -- CP-element group 281: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_req
      -- CP-element group 281: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_992_konst_delay_trans
      -- CP-element group 281: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/$exit
      -- CP-element group 281: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/$exit
      -- 
    phi_stmt_988_req_3424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_988_req_3424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(281), ack => phi_stmt_988_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(281) is a control-delay.
    cp_element_281_delay: control_delay_element  generic map(name => " 281_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(130), ack => convolution3D_CP_1120_elements(281), clk => clk, reset =>reset);
    -- CP-element group 282:  join  transition  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	290 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(280) & convolution3D_CP_1120_elements(281);
      gj_convolution3D_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	138 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (2) 
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Sample/ra
      -- CP-element group 283: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Sample/$exit
      -- 
    ra_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_987_inst_ack_0, ack => convolution3D_CP_1120_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	138 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Update/ca
      -- CP-element group 284: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/Update/$exit
      -- 
    ca_3449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_987_inst_ack_1, ack => convolution3D_CP_1120_elements(284)); -- 
    -- CP-element group 285:  join  transition  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	289 
    -- CP-element group 285:  members (5) 
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_req
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/SplitProtocol/$exit
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/type_cast_987/$exit
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/phi_stmt_981_sources/$exit
      -- CP-element group 285: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_981/$exit
      -- 
    phi_stmt_981_req_3450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_981_req_3450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(285), ack => phi_stmt_981_req_1); -- 
    convolution3D_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(283) & convolution3D_CP_1120_elements(284);
      gj_convolution3D_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	138 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Sample/ra
      -- 
    ra_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_994_inst_ack_0, ack => convolution3D_CP_1120_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	138 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (2) 
      -- CP-element group 287: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/Update/ca
      -- 
    ca_3472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_994_inst_ack_1, ack => convolution3D_CP_1120_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (5) 
      -- CP-element group 288: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/$exit
      -- CP-element group 288: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/$exit
      -- CP-element group 288: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_sources/type_cast_994/SplitProtocol/$exit
      -- CP-element group 288: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/phi_stmt_988_req
      -- CP-element group 288: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_988/$exit
      -- 
    phi_stmt_988_req_3473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_988_req_3473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(288), ack => phi_stmt_988_req_1); -- 
    convolution3D_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(286) & convolution3D_CP_1120_elements(287);
      gj_convolution3D_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	285 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (1) 
      -- CP-element group 289: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(285) & convolution3D_CP_1120_elements(288);
      gj_convolution3D_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  merge  fork  transition  place  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	282 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (2) 
      -- CP-element group 290: 	 branch_block_stmt_436/merge_stmt_980_PhiAck/$entry
      -- CP-element group 290: 	 branch_block_stmt_436/merge_stmt_980_PhiReqMerge
      -- 
    convolution3D_CP_1120_elements(290) <= OrReduce(convolution3D_CP_1120_elements(282) & convolution3D_CP_1120_elements(289));
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (1) 
      -- CP-element group 291: 	 branch_block_stmt_436/merge_stmt_980_PhiAck/phi_stmt_981_ack
      -- 
    phi_stmt_981_ack_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_981_ack_0, ack => convolution3D_CP_1120_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (1) 
      -- CP-element group 292: 	 branch_block_stmt_436/merge_stmt_980_PhiAck/phi_stmt_988_ack
      -- 
    phi_stmt_988_ack_3479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_988_ack_0, ack => convolution3D_CP_1120_elements(292)); -- 
    -- CP-element group 293:  join  fork  transition  place  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	131 
    -- CP-element group 293: 	134 
    -- CP-element group 293: 	135 
    -- CP-element group 293: 	136 
    -- CP-element group 293:  members (16) 
      -- CP-element group 293: 	 branch_block_stmt_436/merge_stmt_980__exit__
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034__entry__
      -- CP-element group 293: 	 branch_block_stmt_436/merge_stmt_980_PhiAck/$exit
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/$entry
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/RPIPE_maxpool_input_pipe_1009_Sample/rr
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_update_start_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1013_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_update_start_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Sample/rr
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1001_to_assign_stmt_1034/type_cast_1028_Update/cr
      -- 
    rr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(293), ack => RPIPE_maxpool_input_pipe_1009_inst_req_0); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(293), ack => type_cast_1013_inst_req_1); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(293), ack => type_cast_1028_inst_req_0); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(293), ack => type_cast_1028_inst_req_1); -- 
    convolution3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(291) & convolution3D_CP_1120_elements(292);
      gj_convolution3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	139 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Sample/ra
      -- CP-element group 294: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Sample/$exit
      -- 
    ra_3503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_0, ack => convolution3D_CP_1120_elements(294)); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	139 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (2) 
      -- CP-element group 295: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/Update/ca
      -- 
    ca_3508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_1, ack => convolution3D_CP_1120_elements(295)); -- 
    -- CP-element group 296:  join  transition  place  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (8) 
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1041_PhiReqMerge
      -- CP-element group 296: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/SplitProtocol/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1045/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/merge_stmt_1041_PhiAck/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1042/phi_stmt_1042_req
      -- 
    phi_stmt_1042_req_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1042_req_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => phi_stmt_1042_req_0); -- 
    convolution3D_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(294) & convolution3D_CP_1120_elements(295);
      gj_convolution3D_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	140 
    -- CP-element group 297: 	141 
    -- CP-element group 297: 	143 
    -- CP-element group 297: 	145 
    -- CP-element group 297:  members (29) 
      -- CP-element group 297: 	 branch_block_stmt_436/merge_stmt_1041__exit__
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080__entry__
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_update_start_
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_resized_1
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_scaled_1
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_computed_1
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_resize_1/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_resize_1/$exit
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_resize_1/index_resize_req
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_resize_1/index_resize_ack
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_scale_1/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_scale_1/$exit
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_scale_1/scale_rename_req
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_index_scale_1/scale_rename_ack
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_update_start
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Sample/req
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/array_obj_ref_1074_final_index_sum_regn_Update/req
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_complete/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/addr_of_1075_complete/req
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_update_start_
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/word_access_complete/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/word_access_complete/word_0/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1052_to_assign_stmt_1080/ptr_deref_1078_Update/word_access_complete/word_0/cr
      -- CP-element group 297: 	 branch_block_stmt_436/merge_stmt_1041_PhiAck/phi_stmt_1042_ack
      -- CP-element group 297: 	 branch_block_stmt_436/merge_stmt_1041_PhiAck/$exit
      -- 
    phi_stmt_1042_ack_3514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1042_ack_0, ack => convolution3D_CP_1120_elements(297)); -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(297), ack => array_obj_ref_1074_index_offset_req_0); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(297), ack => array_obj_ref_1074_index_offset_req_1); -- 
    req_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(297), ack => addr_of_1075_final_reg_req_1); -- 
    cr_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(297), ack => ptr_deref_1078_store_0_req_1); -- 
    -- CP-element group 298:  merge  fork  transition  place  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	129 
    -- CP-element group 298: 	146 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	147 
    -- CP-element group 298: 	148 
    -- CP-element group 298: 	149 
    -- CP-element group 298: 	150 
    -- CP-element group 298: 	151 
    -- CP-element group 298: 	152 
    -- CP-element group 298: 	153 
    -- CP-element group 298: 	154 
    -- CP-element group 298:  members (31) 
      -- CP-element group 298: 	 branch_block_stmt_436/merge_stmt_1082__exit__
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134__entry__
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_update_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1085_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_update_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1089_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_update_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1093_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_update_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1086_to_assign_stmt_1134/type_cast_1097_Update/cr
      -- CP-element group 298: 	 branch_block_stmt_436/merge_stmt_1082_PhiReqMerge
      -- CP-element group 298: 	 branch_block_stmt_436/merge_stmt_1082_PhiAck/dummy
      -- CP-element group 298: 	 branch_block_stmt_436/merge_stmt_1082_PhiAck/$exit
      -- CP-element group 298: 	 branch_block_stmt_436/merge_stmt_1082_PhiAck/$entry
      -- 
    rr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1085_inst_req_0); -- 
    cr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1085_inst_req_1); -- 
    rr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1089_inst_req_0); -- 
    cr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1089_inst_req_1); -- 
    rr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1093_inst_req_0); -- 
    cr_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1093_inst_req_1); -- 
    rr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1097_inst_req_0); -- 
    cr_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => type_cast_1097_inst_req_1); -- 
    convolution3D_CP_1120_elements(298) <= OrReduce(convolution3D_CP_1120_elements(129) & convolution3D_CP_1120_elements(146));
    -- CP-element group 299:  transition  output  delay-element  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	170 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	303 
    -- CP-element group 299:  members (5) 
      -- CP-element group 299: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_req
      -- CP-element group 299: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1219_konst_delay_trans
      -- CP-element group 299: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/$exit
      -- CP-element group 299: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1215/$exit
      -- CP-element group 299: 	 branch_block_stmt_436/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- 
    phi_stmt_1215_req_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1215_req_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(299), ack => phi_stmt_1215_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(299) is a control-delay.
    cp_element_299_delay: control_delay_element  generic map(name => " 299_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(170), ack => convolution3D_CP_1120_elements(299), clk => clk, reset =>reset);
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	212 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Sample/ra
      -- 
    ra_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_0, ack => convolution3D_CP_1120_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	212 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (2) 
      -- CP-element group 301: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/Update/ca
      -- 
    ca_3573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_1, ack => convolution3D_CP_1120_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/SplitProtocol/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_req
      -- CP-element group 302: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/type_cast_1221/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/phi_stmt_1215_sources/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1215/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- 
    phi_stmt_1215_req_3574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1215_req_3574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => phi_stmt_1215_req_1); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(300) & convolution3D_CP_1120_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  merge  transition  place  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	299 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_436/merge_stmt_1214_PhiReqMerge
      -- CP-element group 303: 	 branch_block_stmt_436/merge_stmt_1214_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(303) <= OrReduce(convolution3D_CP_1120_elements(299) & convolution3D_CP_1120_elements(302));
    -- CP-element group 304:  fork  transition  place  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	171 
    -- CP-element group 304: 	172 
    -- CP-element group 304: 	174 
    -- CP-element group 304: 	175 
    -- CP-element group 304: 	178 
    -- CP-element group 304: 	182 
    -- CP-element group 304: 	186 
    -- CP-element group 304: 	190 
    -- CP-element group 304: 	194 
    -- CP-element group 304: 	198 
    -- CP-element group 304: 	202 
    -- CP-element group 304: 	206 
    -- CP-element group 304: 	209 
    -- CP-element group 304:  members (56) 
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_complete/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_resize_1/$exit
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_resize_1/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/addr_of_1228_complete/req
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_computed_1
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Sample/rr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_resize_1/index_resize_req
      -- CP-element group 304: 	 branch_block_stmt_436/merge_stmt_1214__exit__
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377__entry__
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_resize_1/index_resize_ack
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_scale_1/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_scale_1/$exit
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_scale_1/scale_rename_req
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/RPIPE_maxpool_input_pipe_1231_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1248_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_scaled_1
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1320_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Update/req
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1302_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1338_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_final_index_sum_regn_update_start
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1284_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1266_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1235_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_scale_1/scale_rename_ack
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/array_obj_ref_1227_index_resized_1
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/type_cast_1356_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_update_start_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/word_access_complete/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/word_access_complete/word_0/$entry
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1229_to_assign_stmt_1377/ptr_deref_1364_Update/word_access_complete/word_0/cr
      -- CP-element group 304: 	 branch_block_stmt_436/merge_stmt_1214_PhiAck/phi_stmt_1215_ack
      -- CP-element group 304: 	 branch_block_stmt_436/merge_stmt_1214_PhiAck/$exit
      -- 
    phi_stmt_1215_ack_3579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1215_ack_0, ack => convolution3D_CP_1120_elements(304)); -- 
    req_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => addr_of_1228_final_reg_req_1); -- 
    cr_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1248_inst_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1320_inst_req_1); -- 
    cr_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1302_inst_req_1); -- 
    rr_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => RPIPE_maxpool_input_pipe_1231_inst_req_0); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => array_obj_ref_1227_index_offset_req_1); -- 
    cr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1266_inst_req_1); -- 
    cr_2738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1338_inst_req_1); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => array_obj_ref_1227_index_offset_req_0); -- 
    cr_2654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1284_inst_req_1); -- 
    cr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1235_inst_req_1); -- 
    cr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => type_cast_1356_inst_req_1); -- 
    cr_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(304), ack => ptr_deref_1364_store_0_req_1); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	211 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Sample/ra
      -- CP-element group 305: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Sample/$exit
      -- 
    ra_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_0, ack => convolution3D_CP_1120_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	211 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Update/ca
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/Update/$exit
      -- 
    ca_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_1, ack => convolution3D_CP_1120_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_req
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/SplitProtocol/$exit
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1412/$exit
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1409/$exit
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- 
    phi_stmt_1409_req_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1409_req_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(307), ack => phi_stmt_1409_req_0); -- 
    convolution3D_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(305) & convolution3D_CP_1120_elements(306);
      gj_convolution3D_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  transition  output  delay-element  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	157 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (5) 
      -- CP-element group 308: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1409/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_sources/type_cast_1415_konst_delay_trans
      -- CP-element group 308: 	 branch_block_stmt_436/ifx_xend_forx_xend215_PhiReq/phi_stmt_1409/phi_stmt_1409_req
      -- 
    phi_stmt_1409_req_3628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1409_req_3628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(308), ack => phi_stmt_1409_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(308) is a control-delay.
    cp_element_308_delay: control_delay_element  generic map(name => " 308_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(157), ack => convolution3D_CP_1120_elements(308), clk => clk, reset =>reset);
    -- CP-element group 309:  merge  transition  place  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (2) 
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1408_PhiReqMerge
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1408_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(309) <= OrReduce(convolution3D_CP_1120_elements(307) & convolution3D_CP_1120_elements(308));
    -- CP-element group 310:  branch  transition  place  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	213 
    -- CP-element group 310: 	214 
    -- CP-element group 310:  members (15) 
      -- CP-element group 310: 	 branch_block_stmt_436/R_tobool218_1430_place
      -- CP-element group 310: 	 branch_block_stmt_436/merge_stmt_1408__exit__
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1422_to_assign_stmt_1428__entry__
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1422_to_assign_stmt_1428__exit__
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429__entry__
      -- CP-element group 310: 	 branch_block_stmt_436/merge_stmt_1408_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/merge_stmt_1408_PhiAck/phi_stmt_1409_ack
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1422_to_assign_stmt_1428/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1422_to_assign_stmt_1428/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429_dead_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429_eval_test/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429_eval_test/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429_eval_test/branch_req
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429_if_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_436/if_stmt_1429_else_link/$entry
      -- 
    phi_stmt_1409_ack_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1409_ack_0, ack => convolution3D_CP_1120_elements(310)); -- 
    branch_req_2850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(310), ack => if_stmt_1429_branch_req_0); -- 
    -- CP-element group 311:  transition  output  delay-element  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	216 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (4) 
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1458_konst_delay_trans
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_req
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/$exit
      -- 
    phi_stmt_1454_req_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1454_req_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(311), ack => phi_stmt_1454_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(311) is a control-delay.
    cp_element_311_delay: control_delay_element  generic map(name => " 311_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(216), ack => convolution3D_CP_1120_elements(311), clk => clk, reset =>reset);
    -- CP-element group 312:  transition  output  delay-element  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	216 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (4) 
      -- CP-element group 312: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/$exit
      -- CP-element group 312: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$exit
      -- CP-element group 312: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1465_konst_delay_trans
      -- CP-element group 312: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_req
      -- 
    phi_stmt_1461_req_3664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1461_req_3664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(312), ack => phi_stmt_1461_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(312) is a control-delay.
    cp_element_312_delay: control_delay_element  generic map(name => " 312_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(216), ack => convolution3D_CP_1120_elements(312), clk => clk, reset =>reset);
    -- CP-element group 313:  join  transition  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	321 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_436/bbx_xnphx_xi294_forx_xbodyx_xi303_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(311) & convolution3D_CP_1120_elements(312);
      gj_convolution3D_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	224 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Sample/ra
      -- 
    ra_3684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1460_inst_ack_0, ack => convolution3D_CP_1120_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	224 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Update/ca
      -- CP-element group 315: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/Update/$exit
      -- 
    ca_3689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1460_inst_ack_1, ack => convolution3D_CP_1120_elements(315)); -- 
    -- CP-element group 316:  join  transition  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	320 
    -- CP-element group 316:  members (5) 
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/SplitProtocol/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/type_cast_1460/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_sources/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1454/phi_stmt_1454_req
      -- 
    phi_stmt_1454_req_3690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1454_req_3690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(316), ack => phi_stmt_1454_req_1); -- 
    convolution3D_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(314) & convolution3D_CP_1120_elements(315);
      gj_convolution3D_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	224 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/ra
      -- CP-element group 317: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/$exit
      -- 
    ra_3707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_0, ack => convolution3D_CP_1120_elements(317)); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	224 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/ca
      -- 
    ca_3712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_1, ack => convolution3D_CP_1120_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (5) 
      -- CP-element group 319: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_req
      -- CP-element group 319: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/$exit
      -- CP-element group 319: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/$exit
      -- CP-element group 319: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$exit
      -- CP-element group 319: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/phi_stmt_1461/$exit
      -- 
    phi_stmt_1461_req_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1461_req_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(319), ack => phi_stmt_1461_req_1); -- 
    convolution3D_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(317) & convolution3D_CP_1120_elements(318);
      gj_convolution3D_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  transition  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	316 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_436/forx_xbodyx_xi303_forx_xbodyx_xi303_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(316) & convolution3D_CP_1120_elements(319);
      gj_convolution3D_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  merge  fork  transition  place  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	313 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_436/merge_stmt_1453_PhiReqMerge
      -- CP-element group 321: 	 branch_block_stmt_436/merge_stmt_1453_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(321) <= OrReduce(convolution3D_CP_1120_elements(313) & convolution3D_CP_1120_elements(320));
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (1) 
      -- CP-element group 322: 	 branch_block_stmt_436/merge_stmt_1453_PhiAck/phi_stmt_1454_ack
      -- 
    phi_stmt_1454_ack_3718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1454_ack_0, ack => convolution3D_CP_1120_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (1) 
      -- CP-element group 323: 	 branch_block_stmt_436/merge_stmt_1453_PhiAck/phi_stmt_1461_ack
      -- 
    phi_stmt_1461_ack_3719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1461_ack_0, ack => convolution3D_CP_1120_elements(323)); -- 
    -- CP-element group 324:  join  fork  transition  place  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	217 
    -- CP-element group 324: 	220 
    -- CP-element group 324: 	221 
    -- CP-element group 324: 	222 
    -- CP-element group 324:  members (16) 
      -- CP-element group 324: 	 branch_block_stmt_436/merge_stmt_1453__exit__
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507__entry__
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/RPIPE_maxpool_input_pipe_1482_Sample/rr
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_update_start_
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1486_Update/cr
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_update_start_
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Sample/rr
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1474_to_assign_stmt_1507/type_cast_1501_Update/cr
      -- CP-element group 324: 	 branch_block_stmt_436/merge_stmt_1453_PhiAck/$exit
      -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(324), ack => RPIPE_maxpool_input_pipe_1482_inst_req_0); -- 
    cr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(324), ack => type_cast_1486_inst_req_1); -- 
    rr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(324), ack => type_cast_1501_inst_req_0); -- 
    cr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(324), ack => type_cast_1501_inst_req_1); -- 
    convolution3D_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(322) & convolution3D_CP_1120_elements(323);
      gj_convolution3D_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	225 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (2) 
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Sample/ra
      -- CP-element group 325: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Sample/$exit
      -- 
    ra_3743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1518_inst_ack_0, ack => convolution3D_CP_1120_elements(325)); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	225 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (2) 
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/Update/ca
      -- 
    ca_3748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1518_inst_ack_1, ack => convolution3D_CP_1120_elements(326)); -- 
    -- CP-element group 327:  join  transition  place  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (8) 
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1514_PhiReqMerge
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/SplitProtocol/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1518/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/merge_stmt_1514_PhiAck/$entry
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/forx_xbodyx_xi303_getRemainingElementsx_xexit311_PhiReq/$exit
      -- 
    phi_stmt_1515_req_3749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_3749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(327), ack => phi_stmt_1515_req_0); -- 
    convolution3D_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(325) & convolution3D_CP_1120_elements(326);
      gj_convolution3D_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	226 
    -- CP-element group 328: 	227 
    -- CP-element group 328: 	229 
    -- CP-element group 328: 	231 
    -- CP-element group 328:  members (29) 
      -- CP-element group 328: 	 branch_block_stmt_436/merge_stmt_1514__exit__
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553__entry__
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_update_start_
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_resized_1
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_scaled_1
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_computed_1
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_resize_1/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_resize_1/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_resize_1/index_resize_req
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_resize_1/index_resize_ack
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_scale_1/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_scale_1/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_scale_1/scale_rename_req
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_index_scale_1/scale_rename_ack
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_update_start
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Sample/req
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/array_obj_ref_1547_final_index_sum_regn_Update/req
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_complete/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/addr_of_1548_complete/req
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_update_start_
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/word_access_complete/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/word_access_complete/word_0/$entry
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1525_to_assign_stmt_1553/ptr_deref_1551_Update/word_access_complete/word_0/cr
      -- CP-element group 328: 	 branch_block_stmt_436/merge_stmt_1514_PhiAck/phi_stmt_1515_ack
      -- CP-element group 328: 	 branch_block_stmt_436/merge_stmt_1514_PhiAck/$exit
      -- 
    phi_stmt_1515_ack_3754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1515_ack_0, ack => convolution3D_CP_1120_elements(328)); -- 
    req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(328), ack => array_obj_ref_1547_index_offset_req_0); -- 
    req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(328), ack => array_obj_ref_1547_index_offset_req_1); -- 
    req_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(328), ack => addr_of_1548_final_reg_req_1); -- 
    cr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(328), ack => ptr_deref_1551_store_0_req_1); -- 
    -- CP-element group 329:  merge  fork  transition  place  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	213 
    -- CP-element group 329: 	232 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	233 
    -- CP-element group 329: 	234 
    -- CP-element group 329:  members (13) 
      -- CP-element group 329: 	 branch_block_stmt_436/merge_stmt_1555__exit__
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558__entry__
      -- CP-element group 329: 	 branch_block_stmt_436/merge_stmt_1555_PhiReqMerge
      -- CP-element group 329: 	 branch_block_stmt_436/merge_stmt_1555_PhiAck/dummy
      -- CP-element group 329: 	 branch_block_stmt_436/merge_stmt_1555_PhiAck/$exit
      -- CP-element group 329: 	 branch_block_stmt_436/merge_stmt_1555_PhiAck/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_update_start_
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Sample/crr
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/call_stmt_1558/call_stmt_1558_Update/ccr
      -- 
    crr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(329), ack => call_stmt_1558_call_req_0); -- 
    ccr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(329), ack => call_stmt_1558_call_req_1); -- 
    convolution3D_CP_1120_elements(329) <= OrReduce(convolution3D_CP_1120_elements(213) & convolution3D_CP_1120_elements(232));
    -- CP-element group 330:  transition  output  delay-element  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	247 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	334 
    -- CP-element group 330:  members (5) 
      -- CP-element group 330: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1629/$exit
      -- CP-element group 330: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- CP-element group 330: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/$exit
      -- CP-element group 330: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1635_konst_delay_trans
      -- CP-element group 330: 	 branch_block_stmt_436/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_req
      -- 
    phi_stmt_1629_req_3776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1629_req_3776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(330), ack => phi_stmt_1629_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(330) is a control-delay.
    cp_element_330_delay: control_delay_element  generic map(name => " 330_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(247), ack => convolution3D_CP_1120_elements(330), clk => clk, reset =>reset);
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	259 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Sample/ra
      -- 
    ra_3796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1632_inst_ack_0, ack => convolution3D_CP_1120_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	259 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/Update/ca
      -- 
    ca_3801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1632_inst_ack_1, ack => convolution3D_CP_1120_elements(332)); -- 
    -- CP-element group 333:  join  transition  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_sources/type_cast_1632/SplitProtocol/$exit
      -- CP-element group 333: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1629/phi_stmt_1629_req
      -- 
    phi_stmt_1629_req_3802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1629_req_3802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(333), ack => phi_stmt_1629_req_0); -- 
    convolution3D_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(331) & convolution3D_CP_1120_elements(332);
      gj_convolution3D_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  merge  transition  place  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	330 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (2) 
      -- CP-element group 334: 	 branch_block_stmt_436/merge_stmt_1628_PhiReqMerge
      -- CP-element group 334: 	 branch_block_stmt_436/merge_stmt_1628_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(334) <= OrReduce(convolution3D_CP_1120_elements(330) & convolution3D_CP_1120_elements(333));
    -- CP-element group 335:  fork  transition  place  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	248 
    -- CP-element group 335: 	249 
    -- CP-element group 335: 	250 
    -- CP-element group 335: 	251 
    -- CP-element group 335: 	254 
    -- CP-element group 335: 	255 
    -- CP-element group 335: 	256 
    -- CP-element group 335:  members (26) 
      -- CP-element group 335: 	 branch_block_stmt_436/merge_stmt_1628__exit__
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675__entry__
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_update_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1649_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_update_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/type_cast_1653_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_update_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1657_Update/ccr
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_update_start_
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Sample/crr
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1641_to_assign_stmt_1675/call_stmt_1664_Update/ccr
      -- CP-element group 335: 	 branch_block_stmt_436/merge_stmt_1628_PhiAck/$exit
      -- CP-element group 335: 	 branch_block_stmt_436/merge_stmt_1628_PhiAck/phi_stmt_1629_ack
      -- 
    phi_stmt_1629_ack_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1629_ack_0, ack => convolution3D_CP_1120_elements(335)); -- 
    rr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => type_cast_1649_inst_req_0); -- 
    cr_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => type_cast_1649_inst_req_1); -- 
    rr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => type_cast_1653_inst_req_0); -- 
    cr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => type_cast_1653_inst_req_1); -- 
    ccr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => call_stmt_1657_call_req_1); -- 
    crr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => call_stmt_1664_call_req_0); -- 
    ccr_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(335), ack => call_stmt_1664_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1126_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1404_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_935_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1052 : std_logic_vector(63 downto 0);
    signal R_indvar350_1226_resized : std_logic_vector(13 downto 0);
    signal R_indvar350_1226_scaled : std_logic_vector(13 downto 0);
    signal R_indvar364_757_resized : std_logic_vector(13 downto 0);
    signal R_indvar364_757_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1073_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1073_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1546_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1546_scaled : std_logic_vector(13 downto 0);
    signal add102_803 : std_logic_vector(63 downto 0);
    signal add108_821 : std_logic_vector(63 downto 0);
    signal add114_839 : std_logic_vector(63 downto 0);
    signal add120_857 : std_logic_vector(63 downto 0);
    signal add1216x_xi308_1531 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1058 : std_logic_vector(63 downto 0);
    signal add126_875 : std_logic_vector(63 downto 0);
    signal add132_893 : std_logic_vector(63 downto 0);
    signal add13_487 : std_logic_vector(15 downto 0);
    signal add171_1254 : std_logic_vector(63 downto 0);
    signal add177_1272 : std_logic_vector(63 downto 0);
    signal add183_1290 : std_logic_vector(63 downto 0);
    signal add189_1308 : std_logic_vector(63 downto 0);
    signal add195_1326 : std_logic_vector(63 downto 0);
    signal add201_1344 : std_logic_vector(63 downto 0);
    signal add207_1362 : std_logic_vector(63 downto 0);
    signal add23_512 : std_logic_vector(15 downto 0);
    signal add33_537 : std_logic_vector(15 downto 0);
    signal add43_562 : std_logic_vector(15 downto 0);
    signal add53_587 : std_logic_vector(15 downto 0);
    signal add63_612 : std_logic_vector(15 downto 0);
    signal add73_637 : std_logic_vector(15 downto 0);
    signal add96_785 : std_logic_vector(63 downto 0);
    signal add_462 : std_logic_vector(31 downto 0);
    signal addx_xi299_1492 : std_logic_vector(63 downto 0);
    signal addx_xi_1019 : std_logic_vector(63 downto 0);
    signal and217_1422 : std_logic_vector(63 downto 0);
    signal and_953 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1074_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1074_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1074_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1074_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1074_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1074_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1227_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1227_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1227_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1227_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1227_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1227_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_758_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_758_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_758_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_758_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_758_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_758_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1076 : std_logic_vector(31 downto 0);
    signal arrayidx211_1229 : std_logic_vector(31 downto 0);
    signal arrayidx226_1549 : std_logic_vector(31 downto 0);
    signal arrayidx_760 : std_logic_vector(31 downto 0);
    signal call105_812 : std_logic_vector(7 downto 0);
    signal call111_830 : std_logic_vector(7 downto 0);
    signal call117_848 : std_logic_vector(7 downto 0);
    signal call11_478 : std_logic_vector(7 downto 0);
    signal call123_866 : std_logic_vector(7 downto 0);
    signal call129_884 : std_logic_vector(7 downto 0);
    signal call164_1232 : std_logic_vector(7 downto 0);
    signal call168_1245 : std_logic_vector(7 downto 0);
    signal call16_490 : std_logic_vector(7 downto 0);
    signal call174_1263 : std_logic_vector(7 downto 0);
    signal call180_1281 : std_logic_vector(7 downto 0);
    signal call186_1299 : std_logic_vector(7 downto 0);
    signal call192_1317 : std_logic_vector(7 downto 0);
    signal call198_1335 : std_logic_vector(7 downto 0);
    signal call204_1353 : std_logic_vector(7 downto 0);
    signal call21_503 : std_logic_vector(7 downto 0);
    signal call229_1558 : std_logic_vector(63 downto 0);
    signal call26_515 : std_logic_vector(7 downto 0);
    signal call284_1690 : std_logic_vector(63 downto 0);
    signal call2_453 : std_logic_vector(7 downto 0);
    signal call31_528 : std_logic_vector(7 downto 0);
    signal call36_540 : std_logic_vector(7 downto 0);
    signal call41_553 : std_logic_vector(7 downto 0);
    signal call46_565 : std_logic_vector(7 downto 0);
    signal call51_578 : std_logic_vector(7 downto 0);
    signal call56_590 : std_logic_vector(7 downto 0);
    signal call61_603 : std_logic_vector(7 downto 0);
    signal call66_615 : std_logic_vector(7 downto 0);
    signal call6_465 : std_logic_vector(7 downto 0);
    signal call71_628 : std_logic_vector(7 downto 0);
    signal call89_763 : std_logic_vector(7 downto 0);
    signal call93_776 : std_logic_vector(7 downto 0);
    signal call99_794 : std_logic_vector(7 downto 0);
    signal call_440 : std_logic_vector(7 downto 0);
    signal callx_xi297_1483 : std_logic_vector(7 downto 0);
    signal callx_xi_1010 : std_logic_vector(7 downto 0);
    signal cmp161317_1134 : std_logic_vector(0 downto 0);
    signal cmp321_667 : std_logic_vector(0 downto 0);
    signal cmpx_xi302_1507 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1034 : std_logic_vector(0 downto 0);
    signal conv101_798 : std_logic_vector(63 downto 0);
    signal conv107_816 : std_logic_vector(63 downto 0);
    signal conv113_834 : std_logic_vector(63 downto 0);
    signal conv119_852 : std_logic_vector(63 downto 0);
    signal conv125_870 : std_logic_vector(63 downto 0);
    signal conv12_482 : std_logic_vector(15 downto 0);
    signal conv131_888 : std_logic_vector(63 downto 0);
    signal conv145_1086 : std_logic_vector(63 downto 0);
    signal conv147_1090 : std_logic_vector(63 downto 0);
    signal conv150_1094 : std_logic_vector(63 downto 0);
    signal conv153_1098 : std_logic_vector(63 downto 0);
    signal conv155_1128 : std_logic_vector(63 downto 0);
    signal conv165_1236 : std_logic_vector(63 downto 0);
    signal conv170_1249 : std_logic_vector(63 downto 0);
    signal conv176_1267 : std_logic_vector(63 downto 0);
    signal conv182_1285 : std_logic_vector(63 downto 0);
    signal conv188_1303 : std_logic_vector(63 downto 0);
    signal conv194_1321 : std_logic_vector(63 downto 0);
    signal conv19_494 : std_logic_vector(15 downto 0);
    signal conv1_444 : std_logic_vector(31 downto 0);
    signal conv200_1339 : std_logic_vector(63 downto 0);
    signal conv206_1357 : std_logic_vector(63 downto 0);
    signal conv22_507 : std_logic_vector(15 downto 0);
    signal conv230_1687 : std_logic_vector(63 downto 0);
    signal conv255_1650 : std_logic_vector(63 downto 0);
    signal conv261_1654 : std_logic_vector(63 downto 0);
    signal conv285_1695 : std_logic_vector(63 downto 0);
    signal conv29_519 : std_logic_vector(15 downto 0);
    signal conv2x_xi292_1445 : std_logic_vector(31 downto 0);
    signal conv2x_xi_972 : std_logic_vector(31 downto 0);
    signal conv32_532 : std_logic_vector(15 downto 0);
    signal conv39_544 : std_logic_vector(15 downto 0);
    signal conv3_457 : std_logic_vector(31 downto 0);
    signal conv42_557 : std_logic_vector(15 downto 0);
    signal conv49_569 : std_logic_vector(15 downto 0);
    signal conv52_582 : std_logic_vector(15 downto 0);
    signal conv59_594 : std_logic_vector(15 downto 0);
    signal conv5x_xi298_1487 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1014 : std_logic_vector(63 downto 0);
    signal conv62_607 : std_logic_vector(15 downto 0);
    signal conv69_619 : std_logic_vector(15 downto 0);
    signal conv72_632 : std_logic_vector(15 downto 0);
    signal conv79_641 : std_logic_vector(31 downto 0);
    signal conv81_645 : std_logic_vector(31 downto 0);
    signal conv83_661 : std_logic_vector(63 downto 0);
    signal conv90_767 : std_logic_vector(63 downto 0);
    signal conv95_780 : std_logic_vector(63 downto 0);
    signal conv9_469 : std_logic_vector(15 downto 0);
    signal convx_xi301_1502 : std_logic_vector(31 downto 0);
    signal convx_xi_1029 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi296_1461 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_988 : std_logic_vector(63 downto 0);
    signal exitcond32_908 : std_logic_vector(0 downto 0);
    signal exitcond5_1675 : std_logic_vector(0 downto 0);
    signal exitcond_1377 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1007 : std_logic_vector(15 downto 0);
    signal iNsTr_57_1441 : std_logic_vector(63 downto 0);
    signal iNsTr_65_1480 : std_logic_vector(15 downto 0);
    signal iNsTr_73_1525 : std_logic_vector(63 downto 0);
    signal indvar350_1215 : std_logic_vector(63 downto 0);
    signal indvar364_746 : std_logic_vector(63 downto 0);
    signal indvar_1629 : std_logic_vector(31 downto 0);
    signal indvarx_xnext351_1372 : std_logic_vector(63 downto 0);
    signal indvarx_xnext365_903 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1670 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_940 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1409 : std_logic_vector(63 downto 0);
    signal mul148_1103 : std_logic_vector(63 downto 0);
    signal mul151_1108 : std_logic_vector(63 downto 0);
    signal mul154_1113 : std_logic_vector(63 downto 0);
    signal mul236_1564 : std_logic_vector(15 downto 0);
    signal mul249_1569 : std_logic_vector(15 downto 0);
    signal mul254_1641 : std_logic_vector(31 downto 0);
    signal mul260_1646 : std_logic_vector(31 downto 0);
    signal mul82_655 : std_logic_vector(31 downto 0);
    signal mul_650 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi295_1454 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_981 : std_logic_vector(15 downto 0);
    signal phitmp325_1406 : std_logic_vector(63 downto 0);
    signal phitmp_937 : std_logic_vector(63 downto 0);
    signal ptr_deref_1078_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1078_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1078_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1078_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1078_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1078_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1364_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1364_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1364_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1364_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1364_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1364_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1551_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1551_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_895_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_895_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_895_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_895_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_895_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_895_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1119 : std_logic_vector(63 downto 0);
    signal sh_promx_xi309_1537 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1064 : std_logic_vector(63 downto 0);
    signal shl104_809 : std_logic_vector(63 downto 0);
    signal shl10_475 : std_logic_vector(15 downto 0);
    signal shl110_827 : std_logic_vector(63 downto 0);
    signal shl116_845 : std_logic_vector(63 downto 0);
    signal shl122_863 : std_logic_vector(63 downto 0);
    signal shl128_881 : std_logic_vector(63 downto 0);
    signal shl14x_xi310_1542 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1069 : std_logic_vector(63 downto 0);
    signal shl167_1242 : std_logic_vector(63 downto 0);
    signal shl173_1260 : std_logic_vector(63 downto 0);
    signal shl179_1278 : std_logic_vector(63 downto 0);
    signal shl185_1296 : std_logic_vector(63 downto 0);
    signal shl191_1314 : std_logic_vector(63 downto 0);
    signal shl197_1332 : std_logic_vector(63 downto 0);
    signal shl203_1350 : std_logic_vector(63 downto 0);
    signal shl20_500 : std_logic_vector(15 downto 0);
    signal shl30_525 : std_logic_vector(15 downto 0);
    signal shl40_550 : std_logic_vector(15 downto 0);
    signal shl50_575 : std_logic_vector(15 downto 0);
    signal shl60_600 : std_logic_vector(15 downto 0);
    signal shl70_625 : std_logic_vector(15 downto 0);
    signal shl8x_xi300_1498 : std_logic_vector(63 downto 0);
    signal shl8x_xi300x_xlcssa_1515 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1025 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1042 : std_logic_vector(63 downto 0);
    signal shl92_773 : std_logic_vector(63 downto 0);
    signal shl98_791 : std_logic_vector(63 downto 0);
    signal shl_450 : std_logic_vector(31 downto 0);
    signal shlx_xi293_1451 : std_logic_vector(31 downto 0);
    signal shlx_xi_978 : std_logic_vector(31 downto 0);
    signal sub269_1592 : std_logic_vector(15 downto 0);
    signal sub289_1700 : std_logic_vector(63 downto 0);
    signal sub_1586 : std_logic_vector(15 downto 0);
    signal tmp12_1157 : std_logic_vector(63 downto 0);
    signal tmp13_1161 : std_logic_vector(63 downto 0);
    signal tmp14_1166 : std_logic_vector(63 downto 0);
    signal tmp15_1170 : std_logic_vector(63 downto 0);
    signal tmp16_1175 : std_logic_vector(63 downto 0);
    signal tmp17_1179 : std_logic_vector(63 downto 0);
    signal tmp18_1184 : std_logic_vector(63 downto 0);
    signal tmp19_1188 : std_logic_vector(31 downto 0);
    signal tmp20_1193 : std_logic_vector(63 downto 0);
    signal tmp21_1199 : std_logic_vector(63 downto 0);
    signal tmp22_1205 : std_logic_vector(0 downto 0);
    signal tmp24_705 : std_logic_vector(31 downto 0);
    signal tmp25_710 : std_logic_vector(31 downto 0);
    signal tmp26_714 : std_logic_vector(31 downto 0);
    signal tmp27_719 : std_logic_vector(31 downto 0);
    signal tmp28_724 : std_logic_vector(63 downto 0);
    signal tmp29_730 : std_logic_vector(63 downto 0);
    signal tmp30_736 : std_logic_vector(0 downto 0);
    signal tmp326_1474 : std_logic_vector(15 downto 0);
    signal tmp327_1598 : std_logic_vector(15 downto 0);
    signal tmp345_1147 : std_logic_vector(63 downto 0);
    signal tmp346_1153 : std_logic_vector(0 downto 0);
    signal tmp347_1397 : std_logic_vector(63 downto 0);
    signal tmp354_679 : std_logic_vector(31 downto 0);
    signal tmp356_684 : std_logic_vector(31 downto 0);
    signal tmp357_689 : std_logic_vector(63 downto 0);
    signal tmp358_695 : std_logic_vector(63 downto 0);
    signal tmp359_701 : std_logic_vector(0 downto 0);
    signal tmp361_928 : std_logic_vector(63 downto 0);
    signal tmp3_1602 : std_logic_vector(31 downto 0);
    signal tmp4_1608 : std_logic_vector(31 downto 0);
    signal tmp6_1612 : std_logic_vector(31 downto 0);
    signal tmp7_1617 : std_logic_vector(15 downto 0);
    signal tmp8_1621 : std_logic_vector(31 downto 0);
    signal tmp9_1626 : std_logic_vector(31 downto 0);
    signal tmp_1001 : std_logic_vector(15 downto 0);
    signal tobool218_1428 : std_logic_vector(0 downto 0);
    signal tobool_959 : std_logic_vector(0 downto 0);
    signal type_cast_1005_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1023_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1045_wire : std_logic_vector(63 downto 0);
    signal type_cast_1050_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1056_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1062_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1122_wire : std_logic_vector(63 downto 0);
    signal type_cast_1125_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1132_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1145_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1151_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1203_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1210_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1221_wire : std_logic_vector(63 downto 0);
    signal type_cast_1240_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1258_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1294_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1312_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1330_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1348_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1370_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1389_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1395_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1400_wire : std_logic_vector(63 downto 0);
    signal type_cast_1403_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1412_wire : std_logic_vector(63 downto 0);
    signal type_cast_1415_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1426_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1439_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1449_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1458_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1460_wire : std_logic_vector(15 downto 0);
    signal type_cast_1465_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1467_wire : std_logic_vector(63 downto 0);
    signal type_cast_1472_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1478_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1496_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1518_wire : std_logic_vector(63 downto 0);
    signal type_cast_1523_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1529_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1535_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1579_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1584_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1590_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1596_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1606_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1632_wire : std_logic_vector(31 downto 0);
    signal type_cast_1635_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1668_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1685_wire : std_logic_vector(63 downto 0);
    signal type_cast_1693_wire : std_logic_vector(63 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_473_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_498_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_523_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_573_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_598_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_623_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_659_wire : std_logic_vector(63 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_687_wire : std_logic_vector(63 downto 0);
    signal type_cast_693_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_699_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_722_wire : std_logic_vector(63 downto 0);
    signal type_cast_728_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_734_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_741_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_750_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_752_wire : std_logic_vector(63 downto 0);
    signal type_cast_771_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_789_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_807_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_825_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_861_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_879_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_901_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_931_wire : std_logic_vector(63 downto 0);
    signal type_cast_934_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire : std_logic_vector(63 downto 0);
    signal type_cast_946_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_951_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_957_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_970_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_976_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_985_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_987_wire : std_logic_vector(15 downto 0);
    signal type_cast_992_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_994_wire : std_logic_vector(63 downto 0);
    signal type_cast_999_wire_constant : std_logic_vector(15 downto 0);
    signal umax23_1212 : std_logic_vector(63 downto 0);
    signal umax31_743 : std_logic_vector(63 downto 0);
    signal umax360_922 : std_logic_vector(63 downto 0);
    signal umax_1391 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1074_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1074_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1074_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1074_resized_base_address <= "00000000000000";
    array_obj_ref_1227_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1227_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1227_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1227_resized_base_address <= "00000000000000";
    array_obj_ref_1547_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1547_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1547_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1547_resized_base_address <= "00000000000000";
    array_obj_ref_758_constant_part_of_offset <= "00000000000000";
    array_obj_ref_758_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_758_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_758_resized_base_address <= "00000000000000";
    ptr_deref_1078_word_offset_0 <= "00000000000000";
    ptr_deref_1364_word_offset_0 <= "00000000000000";
    ptr_deref_1551_word_offset_0 <= "00000000000000";
    ptr_deref_895_word_offset_0 <= "00000000000000";
    type_cast_1005_wire_constant <= "0000000000000001";
    type_cast_1023_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1050_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1056_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1062_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1117_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1125_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1132_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1145_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1151_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1210_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1240_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1258_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1276_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1294_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1312_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1330_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1348_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1370_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1389_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1395_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1403_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1415_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1426_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1439_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1449_wire_constant <= "00000000000000000000000000000110";
    type_cast_1458_wire_constant <= "0000000000000000";
    type_cast_1465_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1472_wire_constant <= "0000000000000001";
    type_cast_1478_wire_constant <= "0000000000000001";
    type_cast_1496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1523_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1529_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1575_wire_constant <= "11001000";
    type_cast_1579_wire_constant <= "11001000";
    type_cast_1584_wire_constant <= "1111111111111111";
    type_cast_1590_wire_constant <= "1111111111111111";
    type_cast_1596_wire_constant <= "1111111111111111";
    type_cast_1606_wire_constant <= "00000000000000000000000000000001";
    type_cast_1635_wire_constant <= "00000000000000000000000000000000";
    type_cast_1668_wire_constant <= "00000000000000000000000000000001";
    type_cast_448_wire_constant <= "00000000000000000000000000001000";
    type_cast_473_wire_constant <= "0000000000001000";
    type_cast_498_wire_constant <= "0000000000001000";
    type_cast_523_wire_constant <= "0000000000001000";
    type_cast_548_wire_constant <= "0000000000001000";
    type_cast_573_wire_constant <= "0000000000001000";
    type_cast_598_wire_constant <= "0000000000001000";
    type_cast_623_wire_constant <= "0000000000001000";
    type_cast_665_wire_constant <= "00000000000000000000000000000011";
    type_cast_693_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_699_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_728_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_734_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_741_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_750_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_771_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_789_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_807_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_825_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_843_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_861_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_879_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_901_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_934_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_946_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_951_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_957_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_970_wire_constant <= "00000000000000000000000000000001";
    type_cast_976_wire_constant <= "00000000000000000000000000000110";
    type_cast_985_wire_constant <= "0000000000000000";
    type_cast_992_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_999_wire_constant <= "0000000000000001";
    phi_stmt_1042: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1045_wire;
      req(0) <= phi_stmt_1042_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1042",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1042_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1042,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1042
    phi_stmt_1215: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1219_wire_constant & type_cast_1221_wire;
      req <= phi_stmt_1215_req_0 & phi_stmt_1215_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1215",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1215_ack_0,
          idata => idata,
          odata => indvar350_1215,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1215
    phi_stmt_1409: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1412_wire & type_cast_1415_wire_constant;
      req <= phi_stmt_1409_req_0 & phi_stmt_1409_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1409",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1409_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1409,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1409
    phi_stmt_1454: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1458_wire_constant & type_cast_1460_wire;
      req <= phi_stmt_1454_req_0 & phi_stmt_1454_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1454",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1454_ack_0,
          idata => idata,
          odata => nx_x022x_xi295_1454,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1454
    phi_stmt_1461: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1465_wire_constant & type_cast_1467_wire;
      req <= phi_stmt_1461_req_0 & phi_stmt_1461_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1461",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1461_ack_0,
          idata => idata,
          odata => elementx_x021x_xi296_1461,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1461
    phi_stmt_1515: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1518_wire;
      req(0) <= phi_stmt_1515_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1515",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1515_ack_0,
          idata => idata,
          odata => shl8x_xi300x_xlcssa_1515,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1515
    phi_stmt_1629: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1632_wire & type_cast_1635_wire_constant;
      req <= phi_stmt_1629_req_0 & phi_stmt_1629_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1629",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1629_ack_0,
          idata => idata,
          odata => indvar_1629,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1629
    phi_stmt_746: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_750_wire_constant & type_cast_752_wire;
      req <= phi_stmt_746_req_0 & phi_stmt_746_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_746",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_746_ack_0,
          idata => idata,
          odata => indvar364_746,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_746
    phi_stmt_940: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_943_wire & type_cast_946_wire_constant;
      req <= phi_stmt_940_req_0 & phi_stmt_940_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_940",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_940_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_940,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_940
    phi_stmt_981: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_985_wire_constant & type_cast_987_wire;
      req <= phi_stmt_981_req_0 & phi_stmt_981_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_981",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_981_ack_0,
          idata => idata,
          odata => nx_x022x_xi_981,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_981
    phi_stmt_988: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_992_wire_constant & type_cast_994_wire;
      req <= phi_stmt_988_req_0 & phi_stmt_988_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_988",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_988_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_988,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_988
    -- flow-through select operator MUX_1211_inst
    umax23_1212 <= tmp21_1199 when (tmp22_1205(0) /=  '0') else type_cast_1210_wire_constant;
    -- flow-through select operator MUX_1390_inst
    umax_1391 <= tmp345_1147 when (tmp346_1153(0) /=  '0') else type_cast_1389_wire_constant;
    -- flow-through select operator MUX_742_inst
    umax31_743 <= tmp29_730 when (tmp30_736(0) /=  '0') else type_cast_741_wire_constant;
    -- flow-through select operator MUX_921_inst
    umax360_922 <= tmp358_695 when (tmp359_701(0) /=  '0') else type_cast_920_wire_constant;
    addr_of_1075_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1075_final_reg_req_0;
      addr_of_1075_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1075_final_reg_req_1;
      addr_of_1075_final_reg_ack_1<= rack(0);
      addr_of_1075_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1075_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1074_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1076,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1228_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1228_final_reg_req_0;
      addr_of_1228_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1228_final_reg_req_1;
      addr_of_1228_final_reg_ack_1<= rack(0);
      addr_of_1228_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1228_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1227_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1548_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1548_final_reg_req_0;
      addr_of_1548_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1548_final_reg_req_1;
      addr_of_1548_final_reg_ack_1<= rack(0);
      addr_of_1548_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1548_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1547_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_1549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_759_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_759_final_reg_req_0;
      addr_of_759_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_759_final_reg_req_1;
      addr_of_759_final_reg_ack_1<= rack(0);
      addr_of_759_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_759_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_758_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1013_inst_req_0;
      type_cast_1013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1013_inst_req_1;
      type_cast_1013_inst_ack_1<= rack(0);
      type_cast_1013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1014,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1028_inst_req_0;
      type_cast_1028_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1028_inst_req_1;
      type_cast_1028_inst_ack_1<= rack(0);
      type_cast_1028_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1028_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1001,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1029,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1045_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1045_inst_req_0;
      type_cast_1045_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1045_inst_req_1;
      type_cast_1045_inst_ack_1<= rack(0);
      type_cast_1045_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1045_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1025,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1045_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1085_inst_req_0;
      type_cast_1085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1085_inst_req_1;
      type_cast_1085_inst_ack_1<= rack(0);
      type_cast_1085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1089_inst_req_0;
      type_cast_1089_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1089_inst_req_1;
      type_cast_1089_inst_ack_1<= rack(0);
      type_cast_1089_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_637,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1090,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1093_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1093_inst_req_0;
      type_cast_1093_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1093_inst_req_1;
      type_cast_1093_inst_ack_1<= rack(0);
      type_cast_1093_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1093_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_1094,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1097_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1097_inst_req_0;
      type_cast_1097_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1097_inst_req_1;
      type_cast_1097_inst_ack_1<= rack(0);
      type_cast_1097_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1097_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1098,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1122_inst
    process(sext_1119) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1119(63 downto 0);
      type_cast_1122_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1127_inst
    process(ASHR_i64_i64_1126_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1126_wire(63 downto 0);
      conv155_1128 <= tmp_var; -- 
    end process;
    type_cast_1156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1156_inst_req_0;
      type_cast_1156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1156_inst_req_1;
      type_cast_1156_inst_ack_1<= rack(0);
      type_cast_1156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1160_inst_req_0;
      type_cast_1160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1160_inst_req_1;
      type_cast_1160_inst_ack_1<= rack(0);
      type_cast_1160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1169_inst_req_0;
      type_cast_1169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1169_inst_req_1;
      type_cast_1169_inst_ack_1<= rack(0);
      type_cast_1169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1178_inst_req_0;
      type_cast_1178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1178_inst_req_1;
      type_cast_1178_inst_ack_1<= rack(0);
      type_cast_1178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_637,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_1179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1187_inst_req_0;
      type_cast_1187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1187_inst_req_1;
      type_cast_1187_inst_ack_1<= rack(0);
      type_cast_1187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp18_1184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_1188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1192_inst_req_0;
      type_cast_1192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1192_inst_req_1;
      type_cast_1192_inst_ack_1<= rack(0);
      type_cast_1192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1191_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1221_inst_req_0;
      type_cast_1221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1221_inst_req_1;
      type_cast_1221_inst_ack_1<= rack(0);
      type_cast_1221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext351_1372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1221_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1235_inst_req_0;
      type_cast_1235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1235_inst_req_1;
      type_cast_1235_inst_ack_1<= rack(0);
      type_cast_1235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1248_inst_req_0;
      type_cast_1248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1248_inst_req_1;
      type_cast_1248_inst_ack_1<= rack(0);
      type_cast_1248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1266_inst_req_0;
      type_cast_1266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1266_inst_req_1;
      type_cast_1266_inst_ack_1<= rack(0);
      type_cast_1266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1284_inst_req_0;
      type_cast_1284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1284_inst_req_1;
      type_cast_1284_inst_ack_1<= rack(0);
      type_cast_1284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1302_inst_req_0;
      type_cast_1302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1302_inst_req_1;
      type_cast_1302_inst_ack_1<= rack(0);
      type_cast_1302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1338_inst_req_0;
      type_cast_1338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1338_inst_req_1;
      type_cast_1338_inst_ack_1<= rack(0);
      type_cast_1338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1356_inst_req_0;
      type_cast_1356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1356_inst_req_1;
      type_cast_1356_inst_ack_1<= rack(0);
      type_cast_1356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1400_inst
    process(tmp347_1397) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp347_1397(63 downto 0);
      type_cast_1400_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1405_inst
    process(ASHR_i64_i64_1404_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1404_wire(63 downto 0);
      phitmp325_1406 <= tmp_var; -- 
    end process;
    type_cast_1412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1412_inst_req_0;
      type_cast_1412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1412_inst_req_1;
      type_cast_1412_inst_ack_1<= rack(0);
      type_cast_1412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp325_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1412_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1444_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1444_inst_req_0;
      type_cast_1444_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1444_inst_req_1;
      type_cast_1444_inst_ack_1<= rack(0);
      type_cast_1444_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1444_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_57_1441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi292_1445,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1460_inst_req_0;
      type_cast_1460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1460_inst_req_1;
      type_cast_1460_inst_ack_1<= rack(0);
      type_cast_1460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_65_1480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1460_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1467_inst_req_0;
      type_cast_1467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1467_inst_req_1;
      type_cast_1467_inst_ack_1<= rack(0);
      type_cast_1467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi300_1498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1467_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1486_inst_req_0;
      type_cast_1486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1486_inst_req_1;
      type_cast_1486_inst_ack_1<= rack(0);
      type_cast_1486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi297_1483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi298_1487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1501_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1501_inst_req_0;
      type_cast_1501_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1501_inst_req_1;
      type_cast_1501_inst_ack_1<= rack(0);
      type_cast_1501_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1501_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp326_1474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi301_1502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1518_inst_req_0;
      type_cast_1518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1518_inst_req_1;
      type_cast_1518_inst_ack_1<= rack(0);
      type_cast_1518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi300_1498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1518_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1601_inst_req_0;
      type_cast_1601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1601_inst_req_1;
      type_cast_1601_inst_ack_1<= rack(0);
      type_cast_1601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp327_1598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1611_inst_req_0;
      type_cast_1611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1611_inst_req_1;
      type_cast_1611_inst_ack_1<= rack(0);
      type_cast_1611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1620_inst_req_0;
      type_cast_1620_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1620_inst_req_1;
      type_cast_1620_inst_ack_1<= rack(0);
      type_cast_1620_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1620_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1617,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1621,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1632_inst_req_0;
      type_cast_1632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1632_inst_req_1;
      type_cast_1632_inst_ack_1<= rack(0);
      type_cast_1632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1632_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1649_inst_req_0;
      type_cast_1649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1649_inst_req_1;
      type_cast_1649_inst_ack_1<= rack(0);
      type_cast_1649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul254_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1653_inst_req_0;
      type_cast_1653_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1653_inst_req_1;
      type_cast_1653_inst_ack_1<= rack(0);
      type_cast_1653_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1653_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul260_1646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv261_1654,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1686_inst_req_0;
      type_cast_1686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1686_inst_req_1;
      type_cast_1686_inst_ack_1<= rack(0);
      type_cast_1686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1685_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1694_inst_req_0;
      type_cast_1694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1694_inst_req_1;
      type_cast_1694_inst_ack_1<= rack(0);
      type_cast_1694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1693_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv285_1695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_443_inst_req_0;
      type_cast_443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_443_inst_req_1;
      type_cast_443_inst_ack_1<= rack(0);
      type_cast_443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_456_inst_req_0;
      type_cast_456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_456_inst_req_1;
      type_cast_456_inst_ack_1<= rack(0);
      type_cast_456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_468_inst_req_0;
      type_cast_468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_468_inst_req_1;
      type_cast_468_inst_ack_1<= rack(0);
      type_cast_468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_481_inst_req_0;
      type_cast_481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_481_inst_req_1;
      type_cast_481_inst_ack_1<= rack(0);
      type_cast_481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_493_inst_req_0;
      type_cast_493_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_493_inst_req_1;
      type_cast_493_inst_ack_1<= rack(0);
      type_cast_493_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_493_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_490,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_494,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_506_inst_req_0;
      type_cast_506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_506_inst_req_1;
      type_cast_506_inst_ack_1<= rack(0);
      type_cast_506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_507,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_518_inst_req_0;
      type_cast_518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_518_inst_req_1;
      type_cast_518_inst_ack_1<= rack(0);
      type_cast_518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_531_inst_req_0;
      type_cast_531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_531_inst_req_1;
      type_cast_531_inst_ack_1<= rack(0);
      type_cast_531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_543_inst_req_0;
      type_cast_543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_543_inst_req_1;
      type_cast_543_inst_ack_1<= rack(0);
      type_cast_543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_556_inst_req_0;
      type_cast_556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_556_inst_req_1;
      type_cast_556_inst_ack_1<= rack(0);
      type_cast_556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_568_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_568_inst_req_0;
      type_cast_568_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_568_inst_req_1;
      type_cast_568_inst_ack_1<= rack(0);
      type_cast_568_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_568_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_569,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_581_inst_req_0;
      type_cast_581_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_581_inst_req_1;
      type_cast_581_inst_ack_1<= rack(0);
      type_cast_581_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_581_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_578,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_582,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_606_inst_req_0;
      type_cast_606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_606_inst_req_1;
      type_cast_606_inst_ack_1<= rack(0);
      type_cast_606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_618_inst_req_0;
      type_cast_618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_618_inst_req_1;
      type_cast_618_inst_ack_1<= rack(0);
      type_cast_618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_631_inst_req_0;
      type_cast_631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_631_inst_req_1;
      type_cast_631_inst_ack_1<= rack(0);
      type_cast_631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_640_inst_req_0;
      type_cast_640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_640_inst_req_1;
      type_cast_640_inst_ack_1<= rack(0);
      type_cast_640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_644_inst_req_0;
      type_cast_644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_644_inst_req_1;
      type_cast_644_inst_ack_1<= rack(0);
      type_cast_644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_660_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_660_inst_req_0;
      type_cast_660_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_660_inst_req_1;
      type_cast_660_inst_ack_1<= rack(0);
      type_cast_660_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_660_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_659_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_688_inst_req_0;
      type_cast_688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_688_inst_req_1;
      type_cast_688_inst_ack_1<= rack(0);
      type_cast_688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_687_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp357_689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_704_inst_req_0;
      type_cast_704_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_704_inst_req_1;
      type_cast_704_inst_ack_1<= rack(0);
      type_cast_704_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_705,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_713_inst_req_0;
      type_cast_713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_713_inst_req_1;
      type_cast_713_inst_ack_1<= rack(0);
      type_cast_713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp26_714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_723_inst_req_0;
      type_cast_723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_723_inst_req_1;
      type_cast_723_inst_ack_1<= rack(0);
      type_cast_723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_722_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp28_724,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_752_inst_req_0;
      type_cast_752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_752_inst_req_1;
      type_cast_752_inst_ack_1<= rack(0);
      type_cast_752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext365_903,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_752_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_766_inst_req_0;
      type_cast_766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_766_inst_req_1;
      type_cast_766_inst_ack_1<= rack(0);
      type_cast_766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_763,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_779_inst_req_0;
      type_cast_779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_779_inst_req_1;
      type_cast_779_inst_ack_1<= rack(0);
      type_cast_779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_780,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_797_inst_req_0;
      type_cast_797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_797_inst_req_1;
      type_cast_797_inst_ack_1<= rack(0);
      type_cast_797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_794,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_798,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_815_inst_req_0;
      type_cast_815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_815_inst_req_1;
      type_cast_815_inst_ack_1<= rack(0);
      type_cast_815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_833_inst_req_0;
      type_cast_833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_833_inst_req_1;
      type_cast_833_inst_ack_1<= rack(0);
      type_cast_833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_830,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_848,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_869_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_869_inst_req_0;
      type_cast_869_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_869_inst_req_1;
      type_cast_869_inst_ack_1<= rack(0);
      type_cast_869_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_869_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_870,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_931_inst
    process(tmp361_928) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp361_928(63 downto 0);
      type_cast_931_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_936_inst
    process(ASHR_i64_i64_935_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_935_wire(63 downto 0);
      phitmp_937 <= tmp_var; -- 
    end process;
    type_cast_943_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_943_inst_req_0;
      type_cast_943_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_943_inst_req_1;
      type_cast_943_inst_ack_1<= rack(0);
      type_cast_943_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_943_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_937,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_943_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_987_inst_req_0;
      type_cast_987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_987_inst_req_1;
      type_cast_987_inst_ack_1<= rack(0);
      type_cast_987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_987_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1007,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_987_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_994_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_994_inst_req_0;
      type_cast_994_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_994_inst_req_1;
      type_cast_994_inst_ack_1<= rack(0);
      type_cast_994_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_994_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1025,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_994_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1074_index_1_rename
    process(R_ix_x0x_xlcssa_1073_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1073_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1073_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1074_index_1_resize
    process(ix_x0x_xlcssa_940) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_940;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1073_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1074_root_address_inst
    process(array_obj_ref_1074_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1074_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1074_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1227_index_1_rename
    process(R_indvar350_1226_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar350_1226_resized;
      ov(13 downto 0) := iv;
      R_indvar350_1226_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1227_index_1_resize
    process(indvar350_1215) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar350_1215;
      ov := iv(13 downto 0);
      R_indvar350_1226_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1227_root_address_inst
    process(array_obj_ref_1227_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1227_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1227_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1547_index_1_rename
    process(R_ix_x1x_xlcssa_1546_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1546_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1546_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1547_index_1_resize
    process(ix_x1x_xlcssa_1409) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1409;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1546_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1547_root_address_inst
    process(array_obj_ref_1547_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1547_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1547_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_758_index_1_rename
    process(R_indvar364_757_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar364_757_resized;
      ov(13 downto 0) := iv;
      R_indvar364_757_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_758_index_1_resize
    process(indvar364_746) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar364_746;
      ov := iv(13 downto 0);
      R_indvar364_757_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_758_root_address_inst
    process(array_obj_ref_758_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_758_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_758_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1078_addr_0
    process(ptr_deref_1078_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1078_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1078_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1078_base_resize
    process(arrayidx143_1076) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1076;
      ov := iv(13 downto 0);
      ptr_deref_1078_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1078_gather_scatter
    process(shl14x_xi_1069) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1069;
      ov(63 downto 0) := iv;
      ptr_deref_1078_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1078_root_address_inst
    process(ptr_deref_1078_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1078_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1078_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_addr_0
    process(ptr_deref_1364_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1364_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_base_resize
    process(arrayidx211_1229) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1229;
      ov := iv(13 downto 0);
      ptr_deref_1364_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_gather_scatter
    process(add207_1362) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1362;
      ov(63 downto 0) := iv;
      ptr_deref_1364_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1364_root_address_inst
    process(ptr_deref_1364_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1364_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1364_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_addr_0
    process(ptr_deref_1551_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1551_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1551_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_base_resize
    process(arrayidx226_1549) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_1549;
      ov := iv(13 downto 0);
      ptr_deref_1551_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_gather_scatter
    process(shl14x_xi310_1542) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi310_1542;
      ov(63 downto 0) := iv;
      ptr_deref_1551_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_root_address_inst
    process(ptr_deref_1551_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1551_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1551_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_895_addr_0
    process(ptr_deref_895_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_895_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_895_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_895_base_resize
    process(arrayidx_760) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_760;
      ov := iv(13 downto 0);
      ptr_deref_895_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_895_gather_scatter
    process(add132_893) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_893;
      ov(63 downto 0) := iv;
      ptr_deref_895_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_895_root_address_inst
    process(ptr_deref_895_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_895_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_895_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1035_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1034;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1035_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1035_branch_req_0,
          ack0 => if_stmt_1035_branch_ack_0,
          ack1 => if_stmt_1035_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1135_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161317_1134;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1135_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1135_branch_req_0,
          ack0 => if_stmt_1135_branch_ack_0,
          ack1 => if_stmt_1135_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1378_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1377;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1378_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1378_branch_req_0,
          ack0 => if_stmt_1378_branch_ack_0,
          ack1 => if_stmt_1378_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1429_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_1428;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1429_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1429_branch_req_0,
          ack0 => if_stmt_1429_branch_ack_0,
          ack1 => if_stmt_1429_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1508_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi302_1507;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1508_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1508_branch_req_0,
          ack0 => if_stmt_1508_branch_ack_0,
          ack1 => if_stmt_1508_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1676_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1675;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1676_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1676_branch_req_0,
          ack0 => if_stmt_1676_branch_ack_0,
          ack1 => if_stmt_1676_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_668_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp321_667;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_668_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_668_branch_req_0,
          ack0 => if_stmt_668_branch_ack_0,
          ack1 => if_stmt_668_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_909_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond32_908;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_909_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_909_branch_req_0,
          ack0 => if_stmt_909_branch_ack_0,
          ack1 => if_stmt_909_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_960_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_959;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_960_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_960_branch_req_0,
          ack0 => if_stmt_960_branch_ack_0,
          ack1 => if_stmt_960_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1000_inst
    process(nx_x022x_xi_981) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_981, type_cast_999_wire_constant, tmp_var);
      tmp_1001 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1006_inst
    process(nx_x022x_xi_981) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_981, type_cast_1005_wire_constant, tmp_var);
      iNsTr_35_1007 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1473_inst
    process(nx_x022x_xi295_1454) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi295_1454, type_cast_1472_wire_constant, tmp_var);
      tmp326_1474 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1479_inst
    process(nx_x022x_xi295_1454) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi295_1454, type_cast_1478_wire_constant, tmp_var);
      iNsTr_65_1480 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1585_inst
    process(add43_562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43_562, type_cast_1584_wire_constant, tmp_var);
      sub_1586 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1591_inst
    process(add63_612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add63_612, type_cast_1590_wire_constant, tmp_var);
      sub269_1592 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1597_inst
    process(add53_587) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_587, type_cast_1596_wire_constant, tmp_var);
      tmp327_1598 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1607_inst
    process(tmp3_1602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1602, type_cast_1606_wire_constant, tmp_var);
      tmp4_1608 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1645_inst
    process(tmp9_1626, mul254_1641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1626, mul254_1641, tmp_var);
      mul260_1646 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1669_inst
    process(indvar_1629) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1629, type_cast_1668_wire_constant, tmp_var);
      indvarx_xnext_1670 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1371_inst
    process(indvar350_1215) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar350_1215, type_cast_1370_wire_constant, tmp_var);
      indvarx_xnext351_1372 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_902_inst
    process(indvar364_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar364_746, type_cast_901_wire_constant, tmp_var);
      indvarx_xnext365_903 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1450_inst
    process(conv2x_xi292_1445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi292_1445, type_cast_1449_wire_constant, tmp_var);
      shlx_xi293_1451 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_977_inst
    process(conv2x_xi_972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_972, type_cast_976_wire_constant, tmp_var);
      shlx_xi_978 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1057_inst
    process(Bx_xnot_1052) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1052, type_cast_1056_wire_constant, tmp_var);
      add1216x_xi_1058 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1421_inst
    process(conv155_1128) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1128, type_cast_1420_wire_constant, tmp_var);
      and217_1422 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1530_inst
    process(iNsTr_73_1525) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_73_1525, type_cast_1529_wire_constant, tmp_var);
      add1216x_xi308_1531 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_952_inst
    process(conv83_661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_661, type_cast_951_wire_constant, tmp_var);
      and_953 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1126_inst
    process(type_cast_1122_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1122_wire, type_cast_1125_wire_constant, tmp_var);
      ASHR_i64_i64_1126_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1404_inst
    process(type_cast_1400_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1400_wire, type_cast_1403_wire_constant, tmp_var);
      ASHR_i64_i64_1404_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_935_inst
    process(type_cast_931_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_931_wire, type_cast_934_wire_constant, tmp_var);
      ASHR_i64_i64_935_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1674_inst
    process(indvarx_xnext_1670, tmp4_1608) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1670, tmp4_1608, tmp_var);
      exitcond5_1675 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1376_inst
    process(indvarx_xnext351_1372, umax23_1212) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext351_1372, umax23_1212, tmp_var);
      exitcond_1377 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1427_inst
    process(and217_1422) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_1422, type_cast_1426_wire_constant, tmp_var);
      tobool218_1428 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_907_inst
    process(indvarx_xnext365_903, umax31_743) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext365_903, umax31_743, tmp_var);
      exitcond32_908 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_958_inst
    process(and_953) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_953, type_cast_957_wire_constant, tmp_var);
      tobool_959 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1146_inst
    process(conv155_1128) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1128, type_cast_1145_wire_constant, tmp_var);
      tmp345_1147 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1198_inst
    process(tmp20_1193) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1193, type_cast_1197_wire_constant, tmp_var);
      tmp21_1199 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_694_inst
    process(tmp357_689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp357_689, type_cast_693_wire_constant, tmp_var);
      tmp358_695 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_729_inst
    process(tmp28_724) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp28_724, type_cast_728_wire_constant, tmp_var);
      tmp29_730 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1563_inst
    process(add73_637, add23_512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_637, add23_512, tmp_var);
      mul236_1564 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1568_inst
    process(add43_562, add33_537) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add43_562, add33_537, tmp_var);
      mul249_1569 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1616_inst
    process(add73_637, add23_512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_637, add23_512, tmp_var);
      tmp7_1617 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1625_inst
    process(tmp6_1612, tmp8_1621) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1612, tmp8_1621, tmp_var);
      tmp9_1626 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1640_inst
    process(tmp9_1626, indvar_1629) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1626, indvar_1629, tmp_var);
      mul254_1641 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_649_inst
    process(conv79_641, add_462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_641, add_462, tmp_var);
      mul_650 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_654_inst
    process(mul_650, conv81_645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_650, conv81_645, tmp_var);
      mul82_655 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_678_inst
    process(add_462, conv79_641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_462, conv79_641, tmp_var);
      tmp354_679 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_683_inst
    process(tmp354_679, conv81_645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp354_679, conv81_645, tmp_var);
      tmp356_684 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_709_inst
    process(add_462, tmp24_705) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_462, tmp24_705, tmp_var);
      tmp25_710 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_718_inst
    process(tmp25_710, tmp26_714) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_710, tmp26_714, tmp_var);
      tmp27_719 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1102_inst
    process(conv153_1098, conv145_1086) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1098, conv145_1086, tmp_var);
      mul148_1103 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1107_inst
    process(mul148_1103, conv150_1094) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1103, conv150_1094, tmp_var);
      mul151_1108 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1112_inst
    process(mul151_1108, conv147_1090) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1108, conv147_1090, tmp_var);
      mul154_1113 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1165_inst
    process(tmp12_1157, tmp13_1161) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1157, tmp13_1161, tmp_var);
      tmp14_1166 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1174_inst
    process(tmp14_1166, tmp15_1170) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1166, tmp15_1170, tmp_var);
      tmp16_1175 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1183_inst
    process(tmp16_1175, tmp17_1179) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_1175, tmp17_1179, tmp_var);
      tmp18_1184 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_486_inst
    process(shl10_475, conv12_482) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_475, conv12_482, tmp_var);
      add13_487 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_511_inst
    process(shl20_500, conv22_507) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_500, conv22_507, tmp_var);
      add23_512 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_536_inst
    process(shl30_525, conv32_532) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_525, conv32_532, tmp_var);
      add33_537 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_561_inst
    process(shl40_550, conv42_557) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_550, conv42_557, tmp_var);
      add43_562 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_586_inst
    process(shl50_575, conv52_582) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_575, conv52_582, tmp_var);
      add53_587 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_611_inst
    process(shl60_600, conv62_607) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_600, conv62_607, tmp_var);
      add63_612 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_636_inst
    process(shl70_625, conv72_632) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_625, conv72_632, tmp_var);
      add73_637 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_461_inst
    process(shl_450, conv3_457) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_450, conv3_457, tmp_var);
      add_462 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1018_inst
    process(conv5x_xi_1014, elementx_x021x_xi_988) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1014, elementx_x021x_xi_988, tmp_var);
      addx_xi_1019 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1253_inst
    process(shl167_1242, conv170_1249) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1242, conv170_1249, tmp_var);
      add171_1254 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1271_inst
    process(shl173_1260, conv176_1267) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1260, conv176_1267, tmp_var);
      add177_1272 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1289_inst
    process(shl179_1278, conv182_1285) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1278, conv182_1285, tmp_var);
      add183_1290 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1307_inst
    process(shl185_1296, conv188_1303) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1296, conv188_1303, tmp_var);
      add189_1308 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1325_inst
    process(shl191_1314, conv194_1321) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1314, conv194_1321, tmp_var);
      add195_1326 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1343_inst
    process(shl197_1332, conv200_1339) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1332, conv200_1339, tmp_var);
      add201_1344 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1361_inst
    process(shl203_1350, conv206_1357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1350, conv206_1357, tmp_var);
      add207_1362 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1491_inst
    process(conv5x_xi298_1487, elementx_x021x_xi296_1461) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi298_1487, elementx_x021x_xi296_1461, tmp_var);
      addx_xi299_1492 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_784_inst
    process(shl92_773, conv95_780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_773, conv95_780, tmp_var);
      add96_785 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_802_inst
    process(shl98_791, conv101_798) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_791, conv101_798, tmp_var);
      add102_803 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_820_inst
    process(shl104_809, conv107_816) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_809, conv107_816, tmp_var);
      add108_821 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_838_inst
    process(shl110_827, conv113_834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_827, conv113_834, tmp_var);
      add114_839 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_856_inst
    process(shl116_845, conv119_852) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_845, conv119_852, tmp_var);
      add120_857 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_874_inst
    process(shl122_863, conv125_870) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_863, conv125_870, tmp_var);
      add126_875 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_892_inst
    process(shl128_881, conv131_888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_881, conv131_888, tmp_var);
      add132_893 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_474_inst
    process(conv9_469) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_469, type_cast_473_wire_constant, tmp_var);
      shl10_475 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_499_inst
    process(conv19_494) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_494, type_cast_498_wire_constant, tmp_var);
      shl20_500 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_524_inst
    process(conv29_519) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_519, type_cast_523_wire_constant, tmp_var);
      shl30_525 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_549_inst
    process(conv39_544) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_544, type_cast_548_wire_constant, tmp_var);
      shl40_550 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_574_inst
    process(conv49_569) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_569, type_cast_573_wire_constant, tmp_var);
      shl50_575 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_599_inst
    process(conv59_594) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_594, type_cast_598_wire_constant, tmp_var);
      shl60_600 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_624_inst
    process(conv69_619) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_619, type_cast_623_wire_constant, tmp_var);
      shl70_625 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_449_inst
    process(conv1_444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_444, type_cast_448_wire_constant, tmp_var);
      shl_450 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_971_inst
    process(mul82_655) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_655, type_cast_970_wire_constant, tmp_var);
      conv2x_xi_972 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1024_inst
    process(addx_xi_1019) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1019, type_cast_1023_wire_constant, tmp_var);
      shl8x_xi_1025 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1051_inst
    process(conv83_661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_661, type_cast_1050_wire_constant, tmp_var);
      Bx_xnot_1052 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1068_inst
    process(shl8x_xix_xlcssa_1042, sh_promx_xi_1064) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1042, sh_promx_xi_1064, tmp_var);
      shl14x_xi_1069 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1118_inst
    process(mul154_1113) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1113, type_cast_1117_wire_constant, tmp_var);
      sext_1119 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1241_inst
    process(conv165_1236) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1236, type_cast_1240_wire_constant, tmp_var);
      shl167_1242 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1259_inst
    process(add171_1254) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1254, type_cast_1258_wire_constant, tmp_var);
      shl173_1260 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1277_inst
    process(add177_1272) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1272, type_cast_1276_wire_constant, tmp_var);
      shl179_1278 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1295_inst
    process(add183_1290) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1290, type_cast_1294_wire_constant, tmp_var);
      shl185_1296 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1313_inst
    process(add189_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1308, type_cast_1312_wire_constant, tmp_var);
      shl191_1314 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1331_inst
    process(add195_1326) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1326, type_cast_1330_wire_constant, tmp_var);
      shl197_1332 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1349_inst
    process(add201_1344) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1344, type_cast_1348_wire_constant, tmp_var);
      shl203_1350 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1396_inst
    process(umax_1391) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1391, type_cast_1395_wire_constant, tmp_var);
      tmp347_1397 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1440_inst
    process(mul154_1113) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1113, type_cast_1439_wire_constant, tmp_var);
      iNsTr_57_1441 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1497_inst
    process(addx_xi299_1492) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi299_1492, type_cast_1496_wire_constant, tmp_var);
      shl8x_xi300_1498 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1524_inst
    process(mul154_1113) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1113, type_cast_1523_wire_constant, tmp_var);
      iNsTr_73_1525 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1541_inst
    process(shl8x_xi300x_xlcssa_1515, sh_promx_xi309_1537) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi300x_xlcssa_1515, sh_promx_xi309_1537, tmp_var);
      shl14x_xi310_1542 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_772_inst
    process(conv90_767) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_767, type_cast_771_wire_constant, tmp_var);
      shl92_773 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_790_inst
    process(add96_785) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_785, type_cast_789_wire_constant, tmp_var);
      shl98_791 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_808_inst
    process(add102_803) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_803, type_cast_807_wire_constant, tmp_var);
      shl104_809 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_826_inst
    process(add108_821) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_821, type_cast_825_wire_constant, tmp_var);
      shl110_827 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_844_inst
    process(add114_839) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_839, type_cast_843_wire_constant, tmp_var);
      shl116_845 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_862_inst
    process(add120_857) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_857, type_cast_861_wire_constant, tmp_var);
      shl122_863 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_880_inst
    process(add126_875) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_875, type_cast_879_wire_constant, tmp_var);
      shl128_881 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_927_inst
    process(umax360_922) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax360_922, type_cast_926_wire_constant, tmp_var);
      tmp361_928 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1699_inst
    process(conv285_1695, conv230_1687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv285_1695, conv230_1687, tmp_var);
      sub289_1700 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_666_inst
    process(mul82_655) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_655, type_cast_665_wire_constant, tmp_var);
      cmp321_667 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1133_inst
    process(conv155_1128) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1128, type_cast_1132_wire_constant, tmp_var);
      cmp161317_1134 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1152_inst
    process(tmp345_1147) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp345_1147, type_cast_1151_wire_constant, tmp_var);
      tmp346_1153 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1204_inst
    process(tmp21_1199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp21_1199, type_cast_1203_wire_constant, tmp_var);
      tmp22_1205 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_700_inst
    process(tmp358_695) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp358_695, type_cast_699_wire_constant, tmp_var);
      tmp359_701 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_735_inst
    process(tmp29_730) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp29_730, type_cast_734_wire_constant, tmp_var);
      tmp30_736 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1033_inst
    process(convx_xi_1029, shlx_xi_978) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1029, shlx_xi_978, tmp_var);
      cmpx_xi_1034 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1506_inst
    process(convx_xi301_1502, shlx_xi293_1451) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi301_1502, shlx_xi293_1451, tmp_var);
      cmpx_xi302_1507 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1063_inst
    process(add1216x_xi_1058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1058, type_cast_1062_wire_constant, tmp_var);
      sh_promx_xi_1064 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1536_inst
    process(add1216x_xi308_1531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi308_1531, type_cast_1535_wire_constant, tmp_var);
      sh_promx_xi309_1537 <= tmp_var; --
    end process;
    -- shared split operator group (115) : array_obj_ref_1074_index_offset 
    ApIntAdd_group_115: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1073_scaled;
      array_obj_ref_1074_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1074_index_offset_req_0;
      array_obj_ref_1074_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1074_index_offset_req_1;
      array_obj_ref_1074_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_115_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_115_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_115",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 115
    -- shared split operator group (116) : array_obj_ref_1227_index_offset 
    ApIntAdd_group_116: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar350_1226_scaled;
      array_obj_ref_1227_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1227_index_offset_req_0;
      array_obj_ref_1227_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1227_index_offset_req_1;
      array_obj_ref_1227_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_116_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_116_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : array_obj_ref_1547_index_offset 
    ApIntAdd_group_117: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1546_scaled;
      array_obj_ref_1547_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1547_index_offset_req_0;
      array_obj_ref_1547_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1547_index_offset_req_1;
      array_obj_ref_1547_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_117_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : array_obj_ref_758_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar364_757_scaled;
      array_obj_ref_758_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_758_index_offset_req_0;
      array_obj_ref_758_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_758_index_offset_req_1;
      array_obj_ref_758_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- unary operator type_cast_1191_inst
    process(tmp19_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp19_1188, tmp_var);
      type_cast_1191_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1685_inst
    process(call229_1558) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_1558, tmp_var);
      type_cast_1685_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1693_inst
    process(call284_1690) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call284_1690, tmp_var);
      type_cast_1693_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_659_inst
    process(mul82_655) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_655, tmp_var);
      type_cast_659_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_687_inst
    process(tmp356_684) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp356_684, tmp_var);
      type_cast_687_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_722_inst
    process(tmp27_719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp27_719, tmp_var);
      type_cast_722_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_895_store_0 ptr_deref_1078_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_895_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1078_store_0_req_0;
      ptr_deref_895_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1078_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_895_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1078_store_0_req_1;
      ptr_deref_895_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1078_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_895_word_address_0 & ptr_deref_1078_word_address_0;
      data_in <= ptr_deref_895_data_0 & ptr_deref_1078_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1364_store_0 ptr_deref_1551_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1364_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1551_store_0_req_0;
      ptr_deref_1364_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1551_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1364_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1551_store_0_req_1;
      ptr_deref_1364_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1551_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1364_word_address_0 & ptr_deref_1551_word_address_0;
      data_in <= ptr_deref_1364_data_0 & ptr_deref_1551_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_539_inst RPIPE_maxpool_input_pipe_589_inst RPIPE_maxpool_input_pipe_602_inst RPIPE_maxpool_input_pipe_552_inst RPIPE_maxpool_input_pipe_564_inst RPIPE_maxpool_input_pipe_489_inst RPIPE_maxpool_input_pipe_502_inst RPIPE_maxpool_input_pipe_577_inst RPIPE_maxpool_input_pipe_527_inst RPIPE_maxpool_input_pipe_514_inst RPIPE_maxpool_input_pipe_614_inst RPIPE_maxpool_input_pipe_829_inst RPIPE_maxpool_input_pipe_811_inst RPIPE_maxpool_input_pipe_477_inst RPIPE_maxpool_input_pipe_793_inst RPIPE_maxpool_input_pipe_775_inst RPIPE_maxpool_input_pipe_762_inst RPIPE_maxpool_input_pipe_847_inst RPIPE_maxpool_input_pipe_627_inst RPIPE_maxpool_input_pipe_439_inst RPIPE_maxpool_input_pipe_452_inst RPIPE_maxpool_input_pipe_464_inst RPIPE_maxpool_input_pipe_865_inst RPIPE_maxpool_input_pipe_883_inst RPIPE_maxpool_input_pipe_1009_inst RPIPE_maxpool_input_pipe_1231_inst RPIPE_maxpool_input_pipe_1244_inst RPIPE_maxpool_input_pipe_1262_inst RPIPE_maxpool_input_pipe_1280_inst RPIPE_maxpool_input_pipe_1298_inst RPIPE_maxpool_input_pipe_1316_inst RPIPE_maxpool_input_pipe_1334_inst RPIPE_maxpool_input_pipe_1352_inst RPIPE_maxpool_input_pipe_1482_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_539_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_589_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_602_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_552_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_564_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_489_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_502_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_577_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_527_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_514_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_614_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_829_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_811_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_477_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_793_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_775_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_762_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_847_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_627_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_439_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_452_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_464_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_865_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_883_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1009_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1231_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1244_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1262_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1280_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1298_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1316_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1334_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1352_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1482_inst_req_0;
      RPIPE_maxpool_input_pipe_539_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_589_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_602_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_552_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_564_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_489_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_502_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_577_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_527_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_514_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_614_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_829_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_811_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_477_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_793_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_775_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_762_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_847_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_627_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_439_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_452_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_464_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_865_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_883_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1009_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1231_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1244_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1262_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1280_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1298_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1316_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1334_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1352_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1482_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_539_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_589_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_602_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_552_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_564_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_489_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_502_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_577_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_527_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_514_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_614_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_829_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_811_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_477_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_793_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_775_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_762_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_847_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_627_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_439_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_452_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_464_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_865_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_883_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1009_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1231_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1244_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1262_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1280_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1298_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1316_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1334_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1352_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1482_inst_req_1;
      RPIPE_maxpool_input_pipe_539_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_589_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_602_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_552_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_564_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_489_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_502_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_577_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_527_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_514_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_614_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_829_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_811_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_477_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_793_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_775_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_762_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_847_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_627_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_439_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_452_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_464_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_865_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_883_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1009_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1231_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1244_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1262_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1280_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1298_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1316_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1334_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1352_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1482_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call36_540 <= data_out(271 downto 264);
      call56_590 <= data_out(263 downto 256);
      call61_603 <= data_out(255 downto 248);
      call41_553 <= data_out(247 downto 240);
      call46_565 <= data_out(239 downto 232);
      call16_490 <= data_out(231 downto 224);
      call21_503 <= data_out(223 downto 216);
      call51_578 <= data_out(215 downto 208);
      call31_528 <= data_out(207 downto 200);
      call26_515 <= data_out(199 downto 192);
      call66_615 <= data_out(191 downto 184);
      call111_830 <= data_out(183 downto 176);
      call105_812 <= data_out(175 downto 168);
      call11_478 <= data_out(167 downto 160);
      call99_794 <= data_out(159 downto 152);
      call93_776 <= data_out(151 downto 144);
      call89_763 <= data_out(143 downto 136);
      call117_848 <= data_out(135 downto 128);
      call71_628 <= data_out(127 downto 120);
      call_440 <= data_out(119 downto 112);
      call2_453 <= data_out(111 downto 104);
      call6_465 <= data_out(103 downto 96);
      call123_866 <= data_out(95 downto 88);
      call129_884 <= data_out(87 downto 80);
      callx_xi_1010 <= data_out(79 downto 72);
      call164_1232 <= data_out(71 downto 64);
      call168_1245 <= data_out(63 downto 56);
      call174_1263 <= data_out(55 downto 48);
      call180_1281 <= data_out(47 downto 40);
      call186_1299 <= data_out(39 downto 32);
      call192_1317 <= data_out(31 downto 24);
      call198_1335 <= data_out(23 downto 16);
      call204_1353 <= data_out(15 downto 8);
      callx_xi297_1483 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1701_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1701_inst_req_0;
      WPIPE_elapsed_time_pipe_1701_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1701_inst_req_1;
      WPIPE_elapsed_time_pipe_1701_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub289_1700;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_1573_inst WPIPE_maxpool_output_pipe_1577_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1573_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1577_inst_req_0;
      WPIPE_maxpool_output_pipe_1573_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1577_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1573_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1577_inst_req_1;
      WPIPE_maxpool_output_pipe_1573_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1577_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= type_cast_1575_wire_constant & type_cast_1579_wire_constant;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_num_out_pipe_1570_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1570_inst_req_0;
      WPIPE_num_out_pipe_1570_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1570_inst_req_1;
      WPIPE_num_out_pipe_1570_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul249_1569;
      num_out_pipe_write_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_1558_call call_stmt_1690_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1558_call_req_0;
      reqL_unguarded(0) <= call_stmt_1690_call_req_0;
      call_stmt_1558_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1690_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1558_call_req_1;
      reqR_unguarded(0) <= call_stmt_1690_call_req_1;
      call_stmt_1558_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1690_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_1558 <= data_out(127 downto 64);
      call284_1690 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1657_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1657_call_req_0;
      call_stmt_1657_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1657_call_req_1;
      call_stmt_1657_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv255_1650 & conv261_1654;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(127 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1664_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1664_call_req_0;
      call_stmt_1664_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1664_call_req_1;
      call_stmt_1664_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul236_1564 & add33_537 & sub_1586 & sub269_1592 & add23_512 & add13_487;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_3828_start: Boolean;
  signal convolve_CP_3828_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1732_ack_0 : boolean;
  signal nmycount_1791_1731_buf_ack_0 : boolean;
  signal nmycount_1791_1731_buf_req_1 : boolean;
  signal n_out_count_1812_1740_buf_req_0 : boolean;
  signal phi_stmt_1736_req_1 : boolean;
  signal nacc_1783_1735_buf_req_0 : boolean;
  signal n_out_count_1812_1740_buf_req_1 : boolean;
  signal nacc_1783_1735_buf_req_1 : boolean;
  signal n_out_count_1812_1740_buf_ack_0 : boolean;
  signal phi_stmt_1732_req_0 : boolean;
  signal nacc_1783_1735_buf_ack_1 : boolean;
  signal nacc_1783_1735_buf_ack_0 : boolean;
  signal n_out_count_1812_1740_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_1743_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1743_inst_ack_0 : boolean;
  signal phi_stmt_1736_req_0 : boolean;
  signal phi_stmt_1732_req_1 : boolean;
  signal phi_stmt_1736_ack_0 : boolean;
  signal nmycount_1791_1731_buf_req_0 : boolean;
  signal nmycount_1791_1731_buf_ack_1 : boolean;
  signal RPIPE_num_out_pipe_1712_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1712_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1712_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1712_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1715_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1715_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1715_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1715_inst_ack_1 : boolean;
  signal do_while_stmt_1726_branch_req_0 : boolean;
  signal phi_stmt_1728_req_1 : boolean;
  signal phi_stmt_1728_req_0 : boolean;
  signal phi_stmt_1728_ack_0 : boolean;
  signal RPIPE_input_pipe1_1743_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1743_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1750_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1750_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1750_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1750_inst_ack_1 : boolean;
  signal SUB_u32_u32_1764_inst_req_0 : boolean;
  signal SUB_u32_u32_1764_inst_ack_0 : boolean;
  signal SUB_u32_u32_1764_inst_req_1 : boolean;
  signal SUB_u32_u32_1764_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1798_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1798_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1798_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1798_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1819_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_1819_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_1819_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1819_inst_ack_1 : boolean;
  signal slice_1824_inst_req_0 : boolean;
  signal slice_1824_inst_ack_0 : boolean;
  signal slice_1824_inst_req_1 : boolean;
  signal slice_1824_inst_ack_1 : boolean;
  signal slice_1828_inst_req_0 : boolean;
  signal slice_1828_inst_ack_0 : boolean;
  signal slice_1828_inst_req_1 : boolean;
  signal slice_1828_inst_ack_1 : boolean;
  signal W_next_sum_1806_delayed_1_0_1830_inst_req_0 : boolean;
  signal W_next_sum_1806_delayed_1_0_1830_inst_ack_0 : boolean;
  signal W_next_sum_1806_delayed_1_0_1830_inst_req_1 : boolean;
  signal W_next_sum_1806_delayed_1_0_1830_inst_ack_1 : boolean;
  signal type_cast_1836_inst_req_0 : boolean;
  signal type_cast_1836_inst_ack_0 : boolean;
  signal type_cast_1836_inst_req_1 : boolean;
  signal type_cast_1836_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1834_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1834_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1834_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1834_inst_ack_1 : boolean;
  signal W_next_sum_1811_delayed_1_0_1838_inst_req_0 : boolean;
  signal W_next_sum_1811_delayed_1_0_1838_inst_ack_0 : boolean;
  signal W_next_sum_1811_delayed_1_0_1838_inst_req_1 : boolean;
  signal W_next_sum_1811_delayed_1_0_1838_inst_ack_1 : boolean;
  signal type_cast_1844_inst_req_0 : boolean;
  signal type_cast_1844_inst_ack_0 : boolean;
  signal type_cast_1844_inst_req_1 : boolean;
  signal type_cast_1844_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1842_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1842_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1842_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1842_inst_ack_1 : boolean;
  signal do_while_stmt_1726_branch_ack_0 : boolean;
  signal do_while_stmt_1726_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_3828_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3828_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_3828_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3828_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_3828: Block -- control-path 
    signal convolve_CP_3828_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convolve_CP_3828_elements(0) <= convolve_CP_3828_start;
    convolve_CP_3828_symbol <= convolve_CP_3828_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1710/$entry
      -- CP-element group 0: 	 branch_block_stmt_1710/branch_block_stmt_1710__entry__
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725__entry__
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/$entry
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Sample/rr
      -- 
    rr_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(0), ack => RPIPE_num_out_pipe_1712_inst_req_0); -- 
    rr_3864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(0), ack => RPIPE_size_pipe_1715_inst_req_0); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1710/$exit
      -- CP-element group 1: 	 branch_block_stmt_1710/branch_block_stmt_1710__exit__
      -- CP-element group 1: 	 branch_block_stmt_1710/do_while_stmt_1726__exit__
      -- 
    convolve_CP_3828_elements(1) <= convolve_CP_3828_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Update/cr
      -- 
    ra_3851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1712_inst_ack_0, ack => convolve_CP_3828_elements(2)); -- 
    cr_3855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(2), ack => RPIPE_num_out_pipe_1712_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_num_out_pipe_1712_Update/ca
      -- 
    ca_3856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1712_inst_ack_1, ack => convolve_CP_3828_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Update/cr
      -- 
    ra_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1715_inst_ack_0, ack => convolve_CP_3828_elements(4)); -- 
    cr_3869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(4), ack => RPIPE_size_pipe_1715_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/RPIPE_size_pipe_1715_Update/ca
      -- 
    ca_3870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1715_inst_ack_1, ack => convolve_CP_3828_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725__exit__
      -- CP-element group 6: 	 branch_block_stmt_1710/do_while_stmt_1726__entry__
      -- CP-element group 6: 	 branch_block_stmt_1710/assign_stmt_1713_to_assign_stmt_1725/$exit
      -- 
    convolve_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "convolve_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(3) & convolve_CP_3828_elements(5);
      gj_convolve_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1710/do_while_stmt_1726/$entry
      -- CP-element group 7: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726__entry__
      -- 
    convolve_CP_3828_elements(7) <= convolve_CP_3828_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	127 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726__exit__
      -- 
    -- Element group convolve_CP_3828_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_back
      -- 
    -- Element group convolve_CP_3828_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	125 
    -- CP-element group 10: 	126 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1710/do_while_stmt_1726/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_taken/$entry
      -- 
    convolve_CP_3828_elements(10) <= convolve_CP_3828_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	124 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_body_done
      -- 
    convolve_CP_3828_elements(11) <= convolve_CP_3828_elements(124);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	24 
    -- CP-element group 12: 	43 
    -- CP-element group 12: 	62 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_3828_elements(12) <= convolve_CP_3828_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	45 
    -- CP-element group 13: 	64 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_3828_elements(13) <= convolve_CP_3828_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	83 
    -- CP-element group 14: 	123 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_3828_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	123 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/condition_evaluated
      -- 
    condition_evaluated_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(15), ack => do_while_stmt_1726_branch_req_0); -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(19) & convolve_CP_3828_elements(123);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	37 
    -- CP-element group 16: 	56 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	58 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_start__ps
      -- 
    convolve_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(20) & convolve_CP_3828_elements(37) & convolve_CP_3828_elements(56) & convolve_CP_3828_elements(19);
      gj_convolve_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	76 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	84 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	37 
    -- CP-element group 17: 	56 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_completed_
      -- 
    convolve_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(22) & convolve_CP_3828_elements(40) & convolve_CP_3828_elements(59);
      gj_convolve_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	57 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	60 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_start__ps
      -- 
    convolve_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(21) & convolve_CP_3828_elements(38) & convolve_CP_3828_elements(57);
      gj_convolve_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	61 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(23) & convolve_CP_3828_elements(42) & convolve_CP_3828_elements(61);
      gj_convolve_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	86 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_start_
      -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(17) & convolve_CP_3828_elements(86);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	103 
    -- CP-element group 21: 	114 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_start_
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(91) & convolve_CP_3828_elements(103) & convolve_CP_3828_elements(114);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_completed__ps
      -- 
    -- Element group convolve_CP_3828_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	90 
    -- CP-element group 23: 	101 
    -- CP-element group 23: 	112 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_completed__ps
      -- 
    -- Element group convolve_CP_3828_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	12 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_loopback_trigger
      -- 
    convolve_CP_3828_elements(24) <= convolve_CP_3828_elements(12);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_loopback_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_loopback_sample_req_ps
      -- 
    phi_stmt_1728_loopback_sample_req_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_loopback_sample_req_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(25), ack => phi_stmt_1728_req_1); -- 
    -- Element group convolve_CP_3828_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_entry_trigger
      -- 
    convolve_CP_3828_elements(26) <= convolve_CP_3828_elements(13);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_entry_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_entry_sample_req_ps
      -- 
    phi_stmt_1728_entry_sample_req_3903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_entry_sample_req_3903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(27), ack => phi_stmt_1728_req_0); -- 
    -- Element group convolve_CP_3828_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_phi_mux_ack
      -- CP-element group 28: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_phi_mux_ack_ps
      -- 
    phi_stmt_1728_phi_mux_ack_3906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1728_ack_0, ack => convolve_CP_3828_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_sample_completed_
      -- 
    -- Element group convolve_CP_3828_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_update_start_
      -- 
    -- Element group convolve_CP_3828_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_update_completed__ps
      -- 
    convolve_CP_3828_elements(31) <= convolve_CP_3828_elements(32);
    -- CP-element group 32:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	31 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_mcount_var_1730_update_completed_
      -- 
    -- Element group convolve_CP_3828_elements(32) is a control-delay.
    cp_element_32_delay: control_delay_element  generic map(name => " 32_delay", delay_value => 1)  port map(req => convolve_CP_3828_elements(30), ack => convolve_CP_3828_elements(32), clk => clk, reset =>reset);
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_sample_start__ps
      -- 
    req_3927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(33), ack => nmycount_1791_1731_buf_req_0); -- 
    -- Element group convolve_CP_3828_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Update/req
      -- CP-element group 34: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_update_start__ps
      -- 
    req_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(34), ack => nmycount_1791_1731_buf_req_1); -- 
    -- Element group convolve_CP_3828_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Sample/$exit
      -- 
    ack_3928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1791_1731_buf_ack_0, ack => convolve_CP_3828_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nmycount_1731_Update/ack
      -- 
    ack_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1791_1731_buf_ack_1, ack => convolve_CP_3828_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	17 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	16 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_sample_start_
      -- 
    convolve_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(17) & convolve_CP_3828_elements(78) & convolve_CP_3828_elements(82) & convolve_CP_3828_elements(86);
      gj_convolve_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	95 
    -- CP-element group 38: 	99 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	18 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_update_start_
      -- 
    convolve_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(95) & convolve_CP_3828_elements(99);
      gj_convolve_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_sample_start__ps
      -- 
    convolve_CP_3828_elements(39) <= convolve_CP_3828_elements(16);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	17 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_sample_completed__ps
      -- 
    -- Element group convolve_CP_3828_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_update_start__ps
      -- 
    convolve_CP_3828_elements(41) <= convolve_CP_3828_elements(18);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: 	93 
    -- CP-element group 42: 	97 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_update_completed__ps
      -- 
    -- Element group convolve_CP_3828_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	12 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_loopback_trigger
      -- 
    convolve_CP_3828_elements(43) <= convolve_CP_3828_elements(12);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_loopback_sample_req_ps
      -- 
    phi_stmt_1732_loopback_sample_req_3944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1732_loopback_sample_req_3944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(44), ack => phi_stmt_1732_req_1); -- 
    -- Element group convolve_CP_3828_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	13 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_entry_trigger
      -- 
    convolve_CP_3828_elements(45) <= convolve_CP_3828_elements(13);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_entry_sample_req_ps
      -- 
    phi_stmt_1732_entry_sample_req_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1732_entry_sample_req_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(46), ack => phi_stmt_1732_req_0); -- 
    -- Element group convolve_CP_3828_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1732_phi_mux_ack_ps
      -- 
    phi_stmt_1732_phi_mux_ack_3950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1732_ack_0, ack => convolve_CP_3828_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_sample_completed_
      -- 
    -- Element group convolve_CP_3828_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_update_start_
      -- 
    -- Element group convolve_CP_3828_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_update_completed__ps
      -- 
    convolve_CP_3828_elements(50) <= convolve_CP_3828_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_acc_var_1734_update_completed_
      -- 
    -- Element group convolve_CP_3828_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => convolve_CP_3828_elements(49), ack => convolve_CP_3828_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Sample/$entry
      -- 
    req_3971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(52), ack => nacc_1783_1735_buf_req_0); -- 
    -- Element group convolve_CP_3828_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Update/req
      -- CP-element group 53: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_update_start__ps
      -- 
    req_3976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(53), ack => nacc_1783_1735_buf_req_1); -- 
    -- Element group convolve_CP_3828_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_sample_completed__ps
      -- 
    ack_3972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1783_1735_buf_ack_0, ack => convolve_CP_3828_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nacc_1735_update_completed__ps
      -- 
    ack_3977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1783_1735_buf_ack_1, ack => convolve_CP_3828_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	17 
    -- CP-element group 56: 	86 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	16 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_sample_start_
      -- 
    convolve_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(17) & convolve_CP_3828_elements(86);
      gj_convolve_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	88 
    -- CP-element group 57: 	91 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	18 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_update_start_
      -- 
    convolve_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(88) & convolve_CP_3828_elements(91);
      gj_convolve_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_sample_start__ps
      -- 
    convolve_CP_3828_elements(58) <= convolve_CP_3828_elements(16);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_sample_completed__ps
      -- 
    -- Element group convolve_CP_3828_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	18 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_update_start__ps
      -- 
    convolve_CP_3828_elements(60) <= convolve_CP_3828_elements(18);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	87 
    -- CP-element group 61: 	90 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_update_completed__ps
      -- 
    -- Element group convolve_CP_3828_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	12 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_loopback_trigger
      -- 
    convolve_CP_3828_elements(62) <= convolve_CP_3828_elements(12);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_loopback_sample_req_ps
      -- 
    phi_stmt_1736_loopback_sample_req_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1736_loopback_sample_req_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(63), ack => phi_stmt_1736_req_1); -- 
    -- Element group convolve_CP_3828_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	13 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_entry_trigger
      -- 
    convolve_CP_3828_elements(64) <= convolve_CP_3828_elements(13);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_entry_sample_req_ps
      -- CP-element group 65: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_entry_sample_req
      -- 
    phi_stmt_1736_entry_sample_req_3991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1736_entry_sample_req_3991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(65), ack => phi_stmt_1736_req_0); -- 
    -- Element group convolve_CP_3828_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_phi_mux_ack_ps
      -- CP-element group 66: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1736_phi_mux_ack
      -- 
    phi_stmt_1736_phi_mux_ack_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1736_ack_0, ack => convolve_CP_3828_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_sample_start_
      -- 
    -- Element group convolve_CP_3828_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_update_start__ps
      -- 
    -- Element group convolve_CP_3828_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_update_completed__ps
      -- 
    convolve_CP_3828_elements(69) <= convolve_CP_3828_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1739_update_completed_
      -- 
    -- Element group convolve_CP_3828_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convolve_CP_3828_elements(68), ack => convolve_CP_3828_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_sample_start__ps
      -- CP-element group 71: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Sample/$entry
      -- 
    req_4015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(71), ack => n_out_count_1812_1740_buf_req_0); -- 
    -- Element group convolve_CP_3828_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Update/req
      -- CP-element group 72: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_update_start__ps
      -- 
    req_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(72), ack => n_out_count_1812_1740_buf_req_1); -- 
    -- Element group convolve_CP_3828_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_sample_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Sample/$exit
      -- 
    ack_4016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1812_1740_buf_ack_0, ack => convolve_CP_3828_elements(73)); -- 
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_update_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_n_out_count_1740_Update/$exit
      -- 
    ack_4021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1812_1740_buf_ack_1, ack => convolve_CP_3828_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	78 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Sample/rr
      -- 
    rr_4030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(75), ack => RPIPE_input_pipe1_1743_inst_req_0); -- 
    convolve_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(78);
      gj_convolve_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	17 
    -- CP-element group 76: 	77 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	95 
    -- CP-element group 76: 	99 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_update_start_
      -- CP-element group 76: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Update/cr
      -- 
    cr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(76), ack => RPIPE_input_pipe1_1743_inst_req_1); -- 
    convolve_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(17) & convolve_CP_3828_elements(77) & convolve_CP_3828_elements(95) & convolve_CP_3828_elements(99);
      gj_convolve_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	76 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Sample/ra
      -- 
    ra_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1743_inst_ack_0, ack => convolve_CP_3828_elements(77)); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	97 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	75 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_input_pipe1_1743_Update/ca
      -- 
    ca_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1743_inst_ack_1, ack => convolve_CP_3828_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Sample/rr
      -- 
    rr_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(79), ack => RPIPE_kernel_pipe1_1750_inst_req_0); -- 
    convolve_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(82);
      gj_convolve_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: 	81 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	88 
    -- CP-element group 80: 	95 
    -- CP-element group 80: 	99 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_update_start_
      -- CP-element group 80: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Update/cr
      -- 
    cr_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(80), ack => RPIPE_kernel_pipe1_1750_inst_req_1); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(17) & convolve_CP_3828_elements(81) & convolve_CP_3828_elements(88) & convolve_CP_3828_elements(95) & convolve_CP_3828_elements(99);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Sample/ra
      -- 
    ra_4045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1750_inst_ack_0, ack => convolve_CP_3828_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: 	93 
    -- CP-element group 82: 	97 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/RPIPE_kernel_pipe1_1750_Update/ca
      -- 
    ca_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1750_inst_ack_1, ack => convolve_CP_3828_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	14 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Sample/rr
      -- 
    rr_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(83), ack => SUB_u32_u32_1764_inst_req_0); -- 
    convolve_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(14) & convolve_CP_3828_elements(85);
      gj_convolve_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	17 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	103 
    -- CP-element group 84: 	114 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Update/cr
      -- 
    cr_4063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(84), ack => SUB_u32_u32_1764_inst_req_1); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(17) & convolve_CP_3828_elements(91) & convolve_CP_3828_elements(103) & convolve_CP_3828_elements(114);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Sample/ra
      -- 
    ra_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1764_inst_ack_0, ack => convolve_CP_3828_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	90 
    -- CP-element group 86: 	101 
    -- CP-element group 86: 	112 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	20 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	56 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/SUB_u32_u32_1764_Update/ca
      -- 
    ca_4064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1764_inst_ack_1, ack => convolve_CP_3828_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	61 
    -- CP-element group 87: 	82 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Sample/req
      -- 
    req_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(87), ack => WPIPE_kernel_pipe1_1798_inst_req_0); -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(61) & convolve_CP_3828_elements(82) & convolve_CP_3828_elements(89);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	57 
    -- CP-element group 88: 	80 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Sample/ack
      -- CP-element group 88: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Update/req
      -- 
    ack_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1798_inst_ack_0, ack => convolve_CP_3828_elements(88)); -- 
    req_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(88), ack => WPIPE_kernel_pipe1_1798_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	124 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_kernel_pipe1_1798_Update/ack
      -- 
    ack_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1798_inst_ack_1, ack => convolve_CP_3828_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	23 
    -- CP-element group 90: 	61 
    -- CP-element group 90: 	86 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Sample/req
      -- 
    req_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(90), ack => WPIPE_input_done_pipe_1819_inst_req_0); -- 
    convolve_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(23) & convolve_CP_3828_elements(61) & convolve_CP_3828_elements(86) & convolve_CP_3828_elements(92);
      gj_convolve_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	21 
    -- CP-element group 91: 	57 
    -- CP-element group 91: 	84 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Update/req
      -- 
    ack_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1819_inst_ack_0, ack => convolve_CP_3828_elements(91)); -- 
    req_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(91), ack => WPIPE_input_done_pipe_1819_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	124 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_input_done_pipe_1819_Update/ack
      -- 
    ack_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1819_inst_ack_1, ack => convolve_CP_3828_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	42 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	82 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Sample/rr
      -- 
    rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(93), ack => slice_1824_inst_req_0); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(42) & convolve_CP_3828_elements(78) & convolve_CP_3828_elements(82) & convolve_CP_3828_elements(95);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	107 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Update/cr
      -- 
    cr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(94), ack => slice_1824_inst_req_1); -- 
    convolve_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3828_elements(107);
      gj_convolve_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	38 
    -- CP-element group 95: 	76 
    -- CP-element group 95: 	80 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Sample/ra
      -- 
    ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1824_inst_ack_0, ack => convolve_CP_3828_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1824_Update/ca
      -- 
    ca_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1824_inst_ack_1, ack => convolve_CP_3828_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	42 
    -- CP-element group 97: 	78 
    -- CP-element group 97: 	82 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Sample/rr
      -- 
    rr_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(97), ack => slice_1828_inst_req_0); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(42) & convolve_CP_3828_elements(78) & convolve_CP_3828_elements(82) & convolve_CP_3828_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	118 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Update/cr
      -- 
    cr_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(98), ack => slice_1828_inst_req_1); -- 
    convolve_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3828_elements(118);
      gj_convolve_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	38 
    -- CP-element group 99: 	76 
    -- CP-element group 99: 	80 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Sample/ra
      -- 
    ra_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1828_inst_ack_0, ack => convolve_CP_3828_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	116 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/slice_1828_Update/ca
      -- 
    ca_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1828_inst_ack_1, ack => convolve_CP_3828_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	23 
    -- CP-element group 101: 	86 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Sample/req
      -- 
    req_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(101), ack => W_next_sum_1806_delayed_1_0_1830_inst_req_0); -- 
    convolve_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(23) & convolve_CP_3828_elements(86) & convolve_CP_3828_elements(103);
      gj_convolve_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: 	110 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Update/req
      -- 
    req_4133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(102), ack => W_next_sum_1806_delayed_1_0_1830_inst_req_1); -- 
    convolve_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(107) & convolve_CP_3828_elements(110);
      gj_convolve_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	21 
    -- CP-element group 103: 	84 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Sample/ack
      -- 
    ack_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1806_delayed_1_0_1830_inst_ack_0, ack => convolve_CP_3828_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	109 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1832_Update/ack
      -- 
    ack_4134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1806_delayed_1_0_1830_inst_ack_1, ack => convolve_CP_3828_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Sample/rr
      -- 
    rr_4142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(105), ack => type_cast_1836_inst_req_0); -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(96) & convolve_CP_3828_elements(104) & convolve_CP_3828_elements(107);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Update/cr
      -- 
    cr_4147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(106), ack => type_cast_1836_inst_req_1); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3828_elements(110);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Sample/ra
      -- 
    ra_4143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1836_inst_ack_0, ack => convolve_CP_3828_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1836_Update/ca
      -- 
    ca_4148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1836_inst_ack_1, ack => convolve_CP_3828_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	104 
    -- CP-element group 109: 	108 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	122 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Sample/req
      -- 
    req_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(109), ack => WPIPE_maxpool_output_pipe_1834_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(104) & convolve_CP_3828_elements(108) & convolve_CP_3828_elements(122);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	102 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Sample/ack
      -- CP-element group 110: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Update/req
      -- 
    ack_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1834_inst_ack_0, ack => convolve_CP_3828_elements(110)); -- 
    req_4161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(110), ack => WPIPE_maxpool_output_pipe_1834_inst_req_1); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1834_Update/ack
      -- 
    ack_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1834_inst_ack_1, ack => convolve_CP_3828_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	23 
    -- CP-element group 112: 	86 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Sample/req
      -- 
    req_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(112), ack => W_next_sum_1811_delayed_1_0_1838_inst_req_0); -- 
    convolve_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(23) & convolve_CP_3828_elements(86) & convolve_CP_3828_elements(114);
      gj_convolve_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	121 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Update/req
      -- 
    req_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(113), ack => W_next_sum_1811_delayed_1_0_1838_inst_req_1); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(118) & convolve_CP_3828_elements(121);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	21 
    -- CP-element group 114: 	84 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Sample/ack
      -- 
    ack_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1811_delayed_1_0_1838_inst_ack_0, ack => convolve_CP_3828_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/assign_stmt_1840_Update/ack
      -- 
    ack_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1811_delayed_1_0_1838_inst_ack_1, ack => convolve_CP_3828_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	100 
    -- CP-element group 116: 	115 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Sample/rr
      -- 
    rr_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(116), ack => type_cast_1844_inst_req_0); -- 
    convolve_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(100) & convolve_CP_3828_elements(115) & convolve_CP_3828_elements(118);
      gj_convolve_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_update_start_
      -- CP-element group 117: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Update/cr
      -- 
    cr_4189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(117), ack => type_cast_1844_inst_req_1); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_3828_elements(121);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	98 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Sample/ra
      -- 
    ra_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1844_inst_ack_0, ack => convolve_CP_3828_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/type_cast_1844_Update/ca
      -- 
    ca_4190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1844_inst_ack_1, ack => convolve_CP_3828_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Sample/req
      -- 
    req_4198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(120), ack => WPIPE_maxpool_output_pipe_1842_inst_req_0); -- 
    convolve_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(111) & convolve_CP_3828_elements(115) & convolve_CP_3828_elements(119) & convolve_CP_3828_elements(122);
      gj_convolve_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	113 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Update/req
      -- 
    ack_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1842_inst_ack_0, ack => convolve_CP_3828_elements(121)); -- 
    req_4203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3828_elements(121), ack => WPIPE_maxpool_output_pipe_1842_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	109 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/WPIPE_maxpool_output_pipe_1842_Update/ack
      -- 
    ack_4204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1842_inst_ack_1, ack => convolve_CP_3828_elements(122)); -- 
    -- CP-element group 123:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	15 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_3828_elements(123) is a control-delay.
    cp_element_123_delay: control_delay_element  generic map(name => " 123_delay", delay_value => 1)  port map(req => convolve_CP_3828_elements(14), ack => convolve_CP_3828_elements(123), clk => clk, reset =>reset);
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	89 
    -- CP-element group 124: 	92 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	11 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1710/do_while_stmt_1726/do_while_stmt_1726_loop_body/$exit
      -- 
    convolve_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3828_elements(89) & convolve_CP_3828_elements(92) & convolve_CP_3828_elements(122);
      gj_convolve_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3828_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	10 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_exit/$exit
      -- CP-element group 125: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_exit/ack
      -- 
    ack_4209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1726_branch_ack_0, ack => convolve_CP_3828_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	10 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_taken/$exit
      -- CP-element group 126: 	 branch_block_stmt_1710/do_while_stmt_1726/loop_taken/ack
      -- 
    ack_4213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1726_branch_ack_1, ack => convolve_CP_3828_elements(126)); -- 
    -- CP-element group 127:  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1710/do_while_stmt_1726/$exit
      -- 
    convolve_CP_3828_elements(127) <= convolve_CP_3828_elements(8);
    convolve_do_while_stmt_1726_terminator_4214: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1726_terminator_4214", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_3828_elements(11),loop_continue => convolve_CP_3828_elements(126),loop_terminate => convolve_CP_3828_elements(125),loop_back => convolve_CP_3828_elements(9),loop_exit => convolve_CP_3828_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1728_phi_seq_3934_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3828_elements(26);
      convolve_CP_3828_elements(29)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3828_elements(29);
      convolve_CP_3828_elements(30)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3828_elements(31);
      convolve_CP_3828_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3828_elements(24);
      convolve_CP_3828_elements(33)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3828_elements(35);
      convolve_CP_3828_elements(34)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3828_elements(36);
      convolve_CP_3828_elements(25) <= phi_mux_reqs(1);
      phi_stmt_1728_phi_seq_3934 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1728_phi_seq_3934") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3828_elements(16), 
          phi_sample_ack => convolve_CP_3828_elements(22), 
          phi_update_req => convolve_CP_3828_elements(18), 
          phi_update_ack => convolve_CP_3828_elements(23), 
          phi_mux_ack => convolve_CP_3828_elements(28), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1732_phi_seq_3978_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3828_elements(45);
      convolve_CP_3828_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3828_elements(48);
      convolve_CP_3828_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3828_elements(50);
      convolve_CP_3828_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3828_elements(43);
      convolve_CP_3828_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3828_elements(54);
      convolve_CP_3828_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3828_elements(55);
      convolve_CP_3828_elements(44) <= phi_mux_reqs(1);
      phi_stmt_1732_phi_seq_3978 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1732_phi_seq_3978") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3828_elements(39), 
          phi_sample_ack => convolve_CP_3828_elements(40), 
          phi_update_req => convolve_CP_3828_elements(41), 
          phi_update_ack => convolve_CP_3828_elements(42), 
          phi_mux_ack => convolve_CP_3828_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1736_phi_seq_4022_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3828_elements(64);
      convolve_CP_3828_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3828_elements(67);
      convolve_CP_3828_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3828_elements(69);
      convolve_CP_3828_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3828_elements(62);
      convolve_CP_3828_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3828_elements(73);
      convolve_CP_3828_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3828_elements(74);
      convolve_CP_3828_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1736_phi_seq_4022 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1736_phi_seq_4022") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3828_elements(58), 
          phi_sample_ack => convolve_CP_3828_elements(59), 
          phi_update_req => convolve_CP_3828_elements(60), 
          phi_update_ack => convolve_CP_3828_elements(61), 
          phi_mux_ack => convolve_CP_3828_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3886_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_3828_elements(12);
        preds(1)  <= convolve_CP_3828_elements(13);
        entry_tmerge_3886 : transition_merge -- 
          generic map(name => " entry_tmerge_3886")
          port map (preds => preds, symbol_out => convolve_CP_3828_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1808_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_1789_wire : std_logic_vector(31 downto 0);
    signal MUX_1809_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_1744_1744_delayed_1_0_1765 : std_logic_vector(31 downto 0);
    signal acc_1732 : std_logic_vector(15 downto 0);
    signal acc_val_1777 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1829 : std_logic_vector(7 downto 0);
    signal acc_val_up_1825 : std_logic_vector(7 downto 0);
    signal acc_var_1725 : std_logic_vector(15 downto 0);
    signal all_done_flag_1817 : std_logic_vector(0 downto 0);
    signal iread_1744 : std_logic_vector(15 downto 0);
    signal ival_1748 : std_logic_vector(15 downto 0);
    signal konst_1763_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1780_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1786_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1788_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1807_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1820_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1847_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1751 : std_logic_vector(15 downto 0);
    signal kval_1755 : std_logic_vector(15 downto 0);
    signal mcount_var_1720 : std_logic_vector(31 downto 0);
    signal mul_val_1760 : std_logic_vector(15 downto 0);
    signal mycount_1728 : std_logic_vector(31 downto 0);
    signal n_out_count_1812 : std_logic_vector(15 downto 0);
    signal n_out_count_1812_1740_buffered : std_logic_vector(15 downto 0);
    signal nacc_1783 : std_logic_vector(15 downto 0);
    signal nacc_1783_1735_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1770 : std_logic_vector(0 downto 0);
    signal next_sum_1806_delayed_1_0_1832 : std_logic_vector(0 downto 0);
    signal next_sum_1811_delayed_1_0_1840 : std_logic_vector(0 downto 0);
    signal nmycount_1791 : std_logic_vector(31 downto 0);
    signal nmycount_1791_1731_buffered : std_logic_vector(31 downto 0);
    signal num_out_1713 : std_logic_vector(15 downto 0);
    signal out_count_1736 : std_logic_vector(15 downto 0);
    signal out_done_flag_1796 : std_logic_vector(0 downto 0);
    signal size_1716 : std_logic_vector(31 downto 0);
    signal type_cast_1739_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1773_wire : std_logic_vector(15 downto 0);
    signal type_cast_1775_wire : std_logic_vector(15 downto 0);
    signal type_cast_1805_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1836_wire : std_logic_vector(7 downto 0);
    signal type_cast_1844_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1725 <= "0000000000000000";
    konst_1763_wire_constant <= "00000000000000000000000000000001";
    konst_1780_wire_constant <= "0000000000000000";
    konst_1786_wire_constant <= "00000000000000000000000000000000";
    konst_1788_wire_constant <= "00000000000000000000000000000001";
    konst_1807_wire_constant <= "0000000000000001";
    konst_1820_wire_constant <= "1";
    konst_1847_wire_constant <= "1";
    mcount_var_1720 <= "00000000000000000000000000000000";
    type_cast_1739_wire_constant <= "0000000000000001";
    type_cast_1805_wire_constant <= "0000000000000001";
    phi_stmt_1728: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= mcount_var_1720 & nmycount_1791_1731_buffered;
      req <= phi_stmt_1728_req_0 & phi_stmt_1728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1728",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1728_ack_0,
          idata => idata,
          odata => mycount_1728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1728
    phi_stmt_1732: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= acc_var_1725 & nacc_1783_1735_buffered;
      req <= phi_stmt_1732_req_0 & phi_stmt_1732_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1732",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1732_ack_0,
          idata => idata,
          odata => acc_1732,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1732
    phi_stmt_1736: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1739_wire_constant & n_out_count_1812_1740_buffered;
      req <= phi_stmt_1736_req_0 & phi_stmt_1736_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1736",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1736_ack_0,
          idata => idata,
          odata => out_count_1736,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1736
    -- flow-through select operator MUX_1782_inst
    nacc_1783 <= konst_1780_wire_constant when (next_sum_1770(0) /=  '0') else acc_val_1777;
    -- flow-through select operator MUX_1790_inst
    nmycount_1791 <= konst_1786_wire_constant when (next_sum_1770(0) /=  '0') else ADD_u32_u32_1789_wire;
    -- flow-through select operator MUX_1809_inst
    MUX_1809_wire <= type_cast_1805_wire_constant when (out_done_flag_1796(0) /=  '0') else ADD_u16_u16_1808_wire;
    -- flow-through select operator MUX_1811_inst
    n_out_count_1812 <= MUX_1809_wire when (next_sum_1770(0) /=  '0') else out_count_1736;
    slice_1824_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1824_inst_req_0;
      slice_1824_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1824_inst_req_1;
      slice_1824_inst_ack_1<= update_ack(0);
      slice_1824_inst: SliceSplitProtocol generic map(name => "slice_1824_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1777, dout => acc_val_up_1825, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1828_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1828_inst_req_0;
      slice_1828_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1828_inst_req_1;
      slice_1828_inst_ack_1<= update_ack(0);
      slice_1828_inst: SliceSplitProtocol generic map(name => "slice_1828_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1777, dout => acc_val_dn_1829, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1806_delayed_1_0_1830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1806_delayed_1_0_1830_inst_req_0;
      W_next_sum_1806_delayed_1_0_1830_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1806_delayed_1_0_1830_inst_req_1;
      W_next_sum_1806_delayed_1_0_1830_inst_ack_1<= rack(0);
      W_next_sum_1806_delayed_1_0_1830_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1806_delayed_1_0_1830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1806_delayed_1_0_1832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1811_delayed_1_0_1838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1811_delayed_1_0_1838_inst_req_0;
      W_next_sum_1811_delayed_1_0_1838_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1811_delayed_1_0_1838_inst_req_1;
      W_next_sum_1811_delayed_1_0_1838_inst_ack_1<= rack(0);
      W_next_sum_1811_delayed_1_0_1838_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1811_delayed_1_0_1838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1811_delayed_1_0_1840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1812_1740_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1812_1740_buf_req_0;
      n_out_count_1812_1740_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1812_1740_buf_req_1;
      n_out_count_1812_1740_buf_ack_1<= rack(0);
      n_out_count_1812_1740_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1812_1740_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1812_1740_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1783_1735_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1783_1735_buf_req_0;
      nacc_1783_1735_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1783_1735_buf_req_1;
      nacc_1783_1735_buf_ack_1<= rack(0);
      nacc_1783_1735_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1783_1735_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1783_1735_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1791_1731_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1791_1731_buf_req_0;
      nmycount_1791_1731_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1791_1731_buf_req_1;
      nmycount_1791_1731_buf_ack_1<= rack(0);
      nmycount_1791_1731_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1791_1731_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1791_1731_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1747_inst
    process(iread_1744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1744(15 downto 0);
      ival_1748 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1754_inst
    process(kread_1751) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1751(15 downto 0);
      kval_1755 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1773_inst
    process(acc_1732) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1732(15 downto 0);
      type_cast_1773_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1775_inst
    process(mul_val_1760) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1760(15 downto 0);
      type_cast_1775_wire <= tmp_var; -- 
    end process;
    type_cast_1836_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1836_inst_req_0;
      type_cast_1836_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1836_inst_req_1;
      type_cast_1836_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1806_delayed_1_0_1832(0);
      type_cast_1836_inst_gI: SplitGuardInterface generic map(name => "type_cast_1836_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1836_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1836_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1825,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1836_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1844_inst_req_0;
      type_cast_1844_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1844_inst_req_1;
      type_cast_1844_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1811_delayed_1_0_1840(0);
      type_cast_1844_inst_gI: SplitGuardInterface generic map(name => "type_cast_1844_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1844_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1726_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1847_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1726_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1726_branch_req_0,
          ack0 => do_while_stmt_1726_branch_ack_0,
          ack1 => do_while_stmt_1726_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1776_inst
    process(type_cast_1773_wire, type_cast_1775_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1773_wire, type_cast_1775_wire, tmp_var);
      acc_val_1777 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1808_inst
    process(out_count_1736) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1736, konst_1807_wire_constant, tmp_var);
      ADD_u16_u16_1808_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1789_inst
    process(mycount_1728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1728, konst_1788_wire_constant, tmp_var);
      ADD_u32_u32_1789_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1816_inst
    process(out_done_flag_1796, next_sum_1770) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1796, next_sum_1770, tmp_var);
      all_done_flag_1817 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1795_inst
    process(out_count_1736, num_out_1713) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1736, num_out_1713, tmp_var);
      out_done_flag_1796 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1769_inst
    process(mycount_1728, SUB_u32_u32_1744_1744_delayed_1_0_1765) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1728, SUB_u32_u32_1744_1744_delayed_1_0_1765, tmp_var);
      next_sum_1770 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1759_inst
    process(kval_1755, ival_1748) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1755, ival_1748, tmp_var);
      mul_val_1760 <= tmp_var; --
    end process;
    -- shared split operator group (7) : SUB_u32_u32_1764_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1716;
      SUB_u32_u32_1744_1744_delayed_1_0_1765 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_1764_inst_req_0;
      SUB_u32_u32_1764_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_1764_inst_req_1;
      SUB_u32_u32_1764_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared inport operator group (0) : RPIPE_input_pipe1_1743_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1743_inst_req_0;
      RPIPE_input_pipe1_1743_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1743_inst_req_1;
      RPIPE_input_pipe1_1743_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1744 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1750_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1750_inst_req_0;
      RPIPE_kernel_pipe1_1750_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1750_inst_req_1;
      RPIPE_kernel_pipe1_1750_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      kread_1751 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_num_out_pipe_1712_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1712_inst_req_0;
      RPIPE_num_out_pipe_1712_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1712_inst_req_1;
      RPIPE_num_out_pipe_1712_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1713 <= data_out(15 downto 0);
      num_out_pipe_read_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_2: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_size_pipe_1715_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1715_inst_req_0;
      RPIPE_size_pipe_1715_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1715_inst_req_1;
      RPIPE_size_pipe_1715_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_1716 <= data_out(31 downto 0);
      size_pipe_read_3_gI: SplitGuardInterface generic map(name => "size_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_3: InputPortRevised -- 
        generic map ( name => "size_pipe_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1819_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1819_inst_req_0;
      WPIPE_input_done_pipe_1819_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1819_inst_req_1;
      WPIPE_input_done_pipe_1819_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1817(0);
      data_in <= konst_1820_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1798_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1798_inst_req_0;
      WPIPE_kernel_pipe1_1798_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1798_inst_req_1;
      WPIPE_kernel_pipe1_1798_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not out_done_flag_1796(0);
      data_in <= kread_1751;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_maxpool_output_pipe_1834_inst WPIPE_maxpool_output_pipe_1842_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1834_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1842_inst_req_0;
      WPIPE_maxpool_output_pipe_1834_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1842_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1834_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1842_inst_req_1;
      WPIPE_maxpool_output_pipe_1834_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1842_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1811_delayed_1_0_1840(0);
      guard_vector(1)  <= next_sum_1806_delayed_1_0_1832(0);
      data_in <= type_cast_1836_wire & type_cast_1844_wire;
      maxpool_output_pipe_write_2_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_676_start: Boolean;
  signal loadKernelChannel_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nfetch_val_419_358_buf_ack_0 : boolean;
  signal start_add_355_buf_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_1 : boolean;
  signal addr_of_398_final_reg_req_0 : boolean;
  signal addr_of_398_final_reg_ack_0 : boolean;
  signal do_while_stmt_350_branch_ack_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_0 : boolean;
  signal phi_stmt_356_req_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_1 : boolean;
  signal addr_of_398_final_reg_req_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_1 : boolean;
  signal addr_of_398_final_reg_ack_1 : boolean;
  signal type_cast_432_inst_ack_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_0 : boolean;
  signal nfetch_val_419_358_buf_req_0 : boolean;
  signal array_obj_ref_397_index_offset_req_1 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_0 : boolean;
  signal nfetch_val_419_358_buf_req_1 : boolean;
  signal type_cast_432_inst_req_1 : boolean;
  signal do_while_stmt_350_branch_ack_1 : boolean;
  signal my_fetch_339_359_buf_req_1 : boolean;
  signal nfetch_val_419_358_buf_ack_1 : boolean;
  signal my_fetch_339_359_buf_ack_1 : boolean;
  signal my_fetch_339_359_buf_req_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_1 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_0 : boolean;
  signal ptr_deref_406_load_0_ack_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_0 : boolean;
  signal phi_stmt_356_req_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_0 : boolean;
  signal array_obj_ref_397_index_offset_req_0 : boolean;
  signal array_obj_ref_397_index_offset_ack_0 : boolean;
  signal start_add_355_buf_req_1 : boolean;
  signal WPIPE_size_pipe_428_inst_req_1 : boolean;
  signal type_cast_432_inst_req_0 : boolean;
  signal WPIPE_size_pipe_428_inst_req_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_1 : boolean;
  signal array_obj_ref_397_index_offset_ack_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_1 : boolean;
  signal my_fetch_339_359_buf_ack_0 : boolean;
  signal type_cast_432_inst_ack_0 : boolean;
  signal phi_stmt_356_ack_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_0 : boolean;
  signal start_add_355_buf_ack_0 : boolean;
  signal ptr_deref_406_load_0_req_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_1 : boolean;
  signal start_add_355_buf_req_0 : boolean;
  signal array_obj_ref_333_index_offset_req_0 : boolean;
  signal array_obj_ref_333_index_offset_ack_0 : boolean;
  signal array_obj_ref_333_index_offset_req_1 : boolean;
  signal array_obj_ref_333_index_offset_ack_1 : boolean;
  signal addr_of_334_final_reg_req_0 : boolean;
  signal addr_of_334_final_reg_ack_0 : boolean;
  signal addr_of_334_final_reg_req_1 : boolean;
  signal addr_of_334_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_0 : boolean;
  signal ptr_deref_406_load_0_ack_0 : boolean;
  signal ptr_deref_406_load_0_req_0 : boolean;
  signal ptr_deref_338_load_0_req_0 : boolean;
  signal ptr_deref_338_load_0_ack_0 : boolean;
  signal ptr_deref_338_load_0_req_1 : boolean;
  signal ptr_deref_338_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_1 : boolean;
  signal do_while_stmt_350_branch_req_0 : boolean;
  signal phi_stmt_352_req_0 : boolean;
  signal phi_stmt_352_req_1 : boolean;
  signal phi_stmt_352_ack_0 : boolean;
  signal nmycount_374_354_buf_req_0 : boolean;
  signal nmycount_374_354_buf_ack_0 : boolean;
  signal nmycount_374_354_buf_req_1 : boolean;
  signal nmycount_374_354_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_676: Block -- control-path 
    signal loadKernelChannel_CP_676_elements: BooleanArray(94 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_676_elements(0) <= loadKernelChannel_CP_676_start;
    loadKernelChannel_CP_676_symbol <= loadKernelChannel_CP_676_elements(94);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resized_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_computed_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/rr
      -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_0); -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_1); -- 
    cr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => ptr_deref_338_load_0_req_1); -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => RPIPE_input_done_pipe_347_inst_req_0); -- 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => addr_of_334_final_reg_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/ack
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_start_
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_offset_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/req
      -- 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(2)); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(2), ack => addr_of_334_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_completed_
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$exit
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/ack
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_completed_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_start_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_resized
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/rr
      -- 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(4)); -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(4), ack => ptr_deref_338_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_completed_
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/ra
      -- 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_completed_
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_ack
      -- 
    ca_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_completed_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_start_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/ra
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$entry
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/cr
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_0, ack => loadKernelChannel_CP_676_elements(7)); -- 
    cr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(7), ack => RPIPE_input_done_pipe_347_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_completed_
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$exit
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/ca
      -- 
    ca_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_1, ack => loadKernelChannel_CP_676_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_328_to_assign_stmt_348/$exit
      -- CP-element group 9: 	 branch_block_stmt_349/$entry
      -- CP-element group 9: 	 branch_block_stmt_349/branch_block_stmt_349__entry__
      -- CP-element group 9: 	 branch_block_stmt_349/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(8) & loadKernelChannel_CP_676_elements(1) & loadKernelChannel_CP_676_elements(6);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	90 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	91 
    -- CP-element group 10: 	92 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_update_start_
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_sample_start_
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/cr
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/rr
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/$entry
      -- CP-element group 10: 	 assign_stmt_433/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_349/$exit
      -- CP-element group 10: 	 branch_block_stmt_349/branch_block_stmt_349__exit__
      -- CP-element group 10: 	 branch_block_stmt_349/do_while_stmt_350__exit__
      -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_1); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_0); -- 
    loadKernelChannel_CP_676_elements(10) <= loadKernelChannel_CP_676_elements(90);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/$entry
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_CP_676_elements(11) <= loadKernelChannel_CP_676_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	90 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__exit__
      -- 
    -- Element group loadKernelChannel_CP_676_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_349/do_while_stmt_350/loop_back
      -- 
    -- Element group loadKernelChannel_CP_676_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	88 
    -- CP-element group 14: 	89 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/condition_done
      -- 
    loadKernelChannel_CP_676_elements(14) <= loadKernelChannel_CP_676_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	87 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_349/do_while_stmt_350/loop_body_done
      -- 
    loadKernelChannel_CP_676_elements(15) <= loadKernelChannel_CP_676_elements(87);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	47 
    -- CP-element group 16: 	30 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_676_elements(16) <= loadKernelChannel_CP_676_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_676_elements(17) <= loadKernelChannel_CP_676_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	44 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	86 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	29 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/condition_evaluated
      -- 
    condition_evaluated_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(19), ack => do_while_stmt_350_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(86) & loadKernelChannel_CP_676_elements(23) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start__ps
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_req
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(43) & loadKernelChannel_CP_676_elements(24) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	27 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	87 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(45) & loadKernelChannel_CP_676_elements(27);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	44 
    -- CP-element group 22: 	25 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	28 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_req
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(44) & loadKernelChannel_CP_676_elements(25);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	29 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	66 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	80 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(72) & loadKernelChannel_CP_676_elements(80) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start__ps
      -- 
    loadKernelChannel_CP_676_elements(26) <= loadKernelChannel_CP_676_elements(20);
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	21 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start__ps
      -- 
    loadKernelChannel_CP_676_elements(28) <= loadKernelChannel_CP_676_elements(22);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	60 
    -- CP-element group 29: 	66 
    -- CP-element group 29: 	70 
    -- CP-element group 29: 	78 
    -- CP-element group 29: 	19 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (15) 
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed__ps
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(29), ack => array_obj_ref_397_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	16 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(30) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req_ps
      -- 
    phi_stmt_352_loopback_sample_req_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_loopback_sample_req_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(31), ack => phi_stmt_352_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(32) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 33:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req_ps
      -- 
    phi_stmt_352_entry_sample_req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_entry_sample_req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(33), ack => phi_stmt_352_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack_ps
      -- 
    phi_stmt_352_phi_mux_ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_352_ack_0, ack => loadKernelChannel_CP_676_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(35), ack => nmycount_374_354_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start_
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/req
      -- 
    req_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(36), ack => nmycount_374_354_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_0, ack => loadKernelChannel_CP_676_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/ack
      -- 
    ack_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_1, ack => loadKernelChannel_CP_676_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/req
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start__ps
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start_
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(39), ack => start_add_355_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/req
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start__ps
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start_
      -- 
    req_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(40), ack => start_add_355_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed_
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_0, ack => loadKernelChannel_CP_676_elements(41)); -- 
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed__ps
      -- 
    ack_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_1, ack => loadKernelChannel_CP_676_elements(42)); -- 
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	77 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	85 
    -- CP-element group 43: 	21 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start_
      -- 
    loadKernelChannel_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	18 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: 	61 
    -- CP-element group 44: 	84 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	22 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start_
      -- 
    loadKernelChannel_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	21 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	82 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(47) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req
      -- 
    phi_stmt_356_loopback_sample_req_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_loopback_sample_req_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(48), ack => phi_stmt_356_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(49) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req_ps
      -- 
    phi_stmt_356_entry_sample_req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_entry_sample_req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(50), ack => phi_stmt_356_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack_ps
      -- 
    phi_stmt_356_phi_mux_ack_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_356_ack_0, ack => loadKernelChannel_CP_676_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start__ps
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(52), ack => nfetch_val_419_358_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start_
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/req
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start__ps
      -- 
    req_906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(53), ack => nfetch_val_419_358_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed__ps
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_0, ack => loadKernelChannel_CP_676_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed_
      -- 
    ack_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_1, ack => loadKernelChannel_CP_676_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$entry
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(56), ack => my_fetch_339_359_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/req
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start_
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$entry
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(57), ack => my_fetch_339_359_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/ack
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_0, ack => loadKernelChannel_CP_676_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed__ps
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_1, ack => loadKernelChannel_CP_676_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	46 
    -- CP-element group 60: 	29 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$entry
      -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(60), ack => WPIPE_kernel_pipe1_381_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	44 
    -- CP-element group 61: 	25 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_start_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/req
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$exit
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_0, ack => loadKernelChannel_CP_676_elements(61)); -- 
    req_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(61), ack => WPIPE_kernel_pipe1_381_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	87 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$exit
      -- 
    ack_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_1, ack => loadKernelChannel_CP_676_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	67 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$entry
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/req
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_start_
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(63), ack => addr_of_398_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: 	76 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/req
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_start_
      -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(64), ack => addr_of_398_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$entry
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(65), ack => array_obj_ref_397_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	29 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	25 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_sample_complete
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/ack
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (8) 
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_offset_calculated
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_root_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_req
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	65 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$exit
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/ack
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_completed_
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	64 
    -- CP-element group 69:  members (19) 
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_resized
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_calculated
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(70), ack => W_fn_388_delayed_7_0_400_inst_req_0); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(72);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	76 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_start_
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/req
      -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(71), ack => W_fn_388_delayed_7_0_400_inst_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/ack
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_0, ack => loadKernelChannel_CP_676_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/ack
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_1, ack => loadKernelChannel_CP_676_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	73 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$entry
      -- 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(74), ack => ptr_deref_406_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	21 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_start_
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$entry
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(75), ack => ptr_deref_406_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77);
      gj_loadKernelChannel_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	64 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/ra
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$exit
      -- 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	87 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	43 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_ack
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$entry
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$exit
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	29 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/req
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(78), ack => W_fn_394_delayed_13_0_408_inst_req_0); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	21 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/req
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_start_
      -- 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(79), ack => W_fn_394_delayed_13_0_408_inst_req_1); -- 
    loadKernelChannel_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(81);
      gj_loadKernelChannel_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	25 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/ack
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_0, ack => loadKernelChannel_CP_676_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/ack
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$exit
      -- 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_1, ack => loadKernelChannel_CP_676_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	46 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/req
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_start_
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(82), ack => W_fetch_val_396_delayed_13_0_411_inst_req_0); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/req
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_start_
      -- 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(83), ack => W_fetch_val_396_delayed_13_0_411_inst_req_1); -- 
    loadKernelChannel_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	44 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_completed_
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_0, ack => loadKernelChannel_CP_676_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	43 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$exit
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_1, ack => loadKernelChannel_CP_676_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	18 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	19 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_676_elements(18), ack => loadKernelChannel_CP_676_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	62 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	77 
    -- CP-element group 87: 	81 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	21 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(62) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	14 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/ack
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$exit
      -- 
    ack_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_0, ack => loadKernelChannel_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	14 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$exit
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/ack
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_1, ack => loadKernelChannel_CP_676_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	12 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	10 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_349/do_while_stmt_350/$exit
      -- 
    loadKernelChannel_CP_676_elements(90) <= loadKernelChannel_CP_676_elements(12);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	10 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_sample_completed_
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/ra
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_0, ack => loadKernelChannel_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	10 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_start_
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/ca
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/$exit
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/req
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_update_completed_
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$entry
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_1, ack => loadKernelChannel_CP_676_elements(92)); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(92), ack => WPIPE_size_pipe_428_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/ack
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_completed_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_update_start_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/req
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$entry
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$exit
      -- 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_0, ack => loadKernelChannel_CP_676_elements(93)); -- 
    req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(93), ack => WPIPE_size_pipe_428_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/ack
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$exit
      -- CP-element group 94: 	 assign_stmt_433/$exit
      -- CP-element group 94: 	 $exit
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_update_completed_
      -- 
    ack_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_1, ack => loadKernelChannel_CP_676_elements(94)); -- 
    loadKernelChannel_do_while_stmt_350_terminator_1088: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_350_terminator_1088", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_676_elements(15),loop_continue => loadKernelChannel_CP_676_elements(89),loop_terminate => loadKernelChannel_CP_676_elements(88),loop_back => loadKernelChannel_CP_676_elements(13),loop_exit => loadKernelChannel_CP_676_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_352_phi_seq_872_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(30);
      loadKernelChannel_CP_676_elements(35)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(37);
      loadKernelChannel_CP_676_elements(36)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(38);
      loadKernelChannel_CP_676_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(32);
      loadKernelChannel_CP_676_elements(39)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(41);
      loadKernelChannel_CP_676_elements(40)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(42);
      loadKernelChannel_CP_676_elements(33) <= phi_mux_reqs(1);
      phi_stmt_352_phi_seq_872 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_352_phi_seq_872") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(26), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(27), 
          phi_update_req => loadKernelChannel_CP_676_elements(28), 
          phi_update_ack => loadKernelChannel_CP_676_elements(29), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(34), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_356_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(47);
      loadKernelChannel_CP_676_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(54);
      loadKernelChannel_CP_676_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(55);
      loadKernelChannel_CP_676_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(49);
      loadKernelChannel_CP_676_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(58);
      loadKernelChannel_CP_676_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(59);
      loadKernelChannel_CP_676_elements(50) <= phi_mux_reqs(1);
      phi_stmt_356_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_356_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(45), 
          phi_update_req => loadKernelChannel_CP_676_elements(22), 
          phi_update_ack => loadKernelChannel_CP_676_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_814_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_676_elements(16);
        preds(1)  <= loadKernelChannel_CP_676_elements(17);
        entry_tmerge_814 : transition_merge -- 
          generic map(name => " entry_tmerge_814")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_676_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_365_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_387_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_378_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_396_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_332_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_332_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_366_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_424_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_431_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_425_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_333_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_335 : std_logic_vector(31 downto 0);
    signal fetch_addr_399 : std_logic_vector(31 downto 0);
    signal fetch_val_356 : std_logic_vector(63 downto 0);
    signal fetch_val_396_delayed_13_0_413 : std_logic_vector(63 downto 0);
    signal first_fill_344 : std_logic_vector(0 downto 0);
    signal fn_388_delayed_7_0_402 : std_logic_vector(0 downto 0);
    signal fn_390 : std_logic_vector(0 downto 0);
    signal fn_394_delayed_13_0_410 : std_logic_vector(0 downto 0);
    signal fv_407 : std_logic_vector(63 downto 0);
    signal konst_326_wire_constant : std_logic_vector(63 downto 0);
    signal konst_342_wire_constant : std_logic_vector(63 downto 0);
    signal konst_362_wire_constant : std_logic_vector(63 downto 0);
    signal konst_364_wire_constant : std_logic_vector(63 downto 0);
    signal konst_367_wire_constant : std_logic_vector(63 downto 0);
    signal konst_372_wire_constant : std_logic_vector(63 downto 0);
    signal konst_386_wire_constant : std_logic_vector(63 downto 0);
    signal konst_388_wire_constant : std_logic_vector(63 downto 0);
    signal konst_395_wire_constant : std_logic_vector(63 downto 0);
    signal konst_423_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_339 : std_logic_vector(63 downto 0);
    signal my_fetch_339_359_buffered : std_logic_vector(63 downto 0);
    signal my_num1_369 : std_logic_vector(63 downto 0);
    signal mycount_352 : std_logic_vector(63 downto 0);
    signal nfetch_val_419 : std_logic_vector(63 downto 0);
    signal nfetch_val_419_358_buffered : std_logic_vector(63 downto 0);
    signal nmycount_374 : std_logic_vector(63 downto 0);
    signal nmycount_374_354_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_338_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_338_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_406_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_328 : std_logic_vector(63 downto 0);
    signal start_add_355_buffered : std_logic_vector(63 downto 0);
    signal start_next_348 : std_logic_vector(0 downto 0);
    signal type_cast_432_wire : std_logic_vector(31 downto 0);
    signal var_val_380 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_333_constant_part_of_offset <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_333_resized_base_address <= "00000000000000";
    array_obj_ref_397_constant_part_of_offset <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_397_resized_base_address <= "00000000000000";
    konst_326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_367_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_395_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_338_word_offset_0 <= "00000000000000";
    ptr_deref_406_word_offset_0 <= "00000000000000";
    phi_stmt_352: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_374_354_buffered & start_add_355_buffered;
      req <= phi_stmt_352_req_0 & phi_stmt_352_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_352",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_352_ack_0,
          idata => idata,
          odata => mycount_352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_352
    phi_stmt_356: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_419_358_buffered & my_fetch_339_359_buffered;
      req <= phi_stmt_356_req_0 & phi_stmt_356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_356",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_356_ack_0,
          idata => idata,
          odata => fetch_val_356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_356
    -- flow-through select operator MUX_418_inst
    nfetch_val_419 <= fv_407 when (fn_394_delayed_13_0_410(0) /=  '0') else fetch_val_396_delayed_13_0_413;
    W_fetch_val_396_delayed_13_0_411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_0;
      W_fetch_val_396_delayed_13_0_411_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_1;
      W_fetch_val_396_delayed_13_0_411_inst_ack_1<= rack(0);
      W_fetch_val_396_delayed_13_0_411_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_396_delayed_13_0_411_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_396_delayed_13_0_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_388_delayed_7_0_400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_388_delayed_7_0_400_inst_req_0;
      W_fn_388_delayed_7_0_400_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_388_delayed_7_0_400_inst_req_1;
      W_fn_388_delayed_7_0_400_inst_ack_1<= rack(0);
      W_fn_388_delayed_7_0_400_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_388_delayed_7_0_400_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_388_delayed_7_0_402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_394_delayed_13_0_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_394_delayed_13_0_408_inst_req_0;
      W_fn_394_delayed_13_0_408_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_394_delayed_13_0_408_inst_req_1;
      W_fn_394_delayed_13_0_408_inst_ack_1<= rack(0);
      W_fn_394_delayed_13_0_408_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_394_delayed_13_0_408_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_394_delayed_13_0_410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_334_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_334_final_reg_req_0;
      addr_of_334_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_334_final_reg_req_1;
      addr_of_334_final_reg_ack_1<= rack(0);
      addr_of_334_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_334_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_333_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_398_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_398_final_reg_req_0;
      addr_of_398_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_398_final_reg_req_1;
      addr_of_398_final_reg_ack_1<= rack(0);
      addr_of_398_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_398_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_397_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_339_359_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_339_359_buf_req_0;
      my_fetch_339_359_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_339_359_buf_req_1;
      my_fetch_339_359_buf_ack_1<= rack(0);
      my_fetch_339_359_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_339_359_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_339_359_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_419_358_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_419_358_buf_req_0;
      nfetch_val_419_358_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_419_358_buf_req_1;
      nfetch_val_419_358_buf_ack_1<= rack(0);
      nfetch_val_419_358_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_419_358_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_419_358_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_374_354_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_374_354_buf_req_0;
      nmycount_374_354_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_374_354_buf_req_1;
      nmycount_374_354_buf_ack_1<= rack(0);
      nmycount_374_354_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_374_354_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_374_354_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_355_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_355_buf_req_0;
      start_add_355_buf_ack_0<= wack(0);
      rreq(0) <= start_add_355_buf_req_1;
      start_add_355_buf_ack_1<= rack(0);
      start_add_355_buf : InterlockBuffer generic map ( -- 
        name => "start_add_355_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_355_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_379_inst
    process(LSHR_u64_u64_378_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_378_wire(15 downto 0);
      var_val_380 <= tmp_var; -- 
    end process;
    type_cast_432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_432_inst_req_0;
      type_cast_432_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_432_inst_req_1;
      type_cast_432_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  first_fill_344(0);
      type_cast_432_inst_gI: SplitGuardInterface generic map(name => "type_cast_432_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SUB_u64_u64_431_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_333_index_1_rename
    process(R_sh_start_332_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_332_resized;
      ov(13 downto 0) := iv;
      R_sh_start_332_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_index_1_resize
    process(sh_start_328) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_328;
      ov := iv(13 downto 0);
      R_sh_start_332_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_root_address_inst
    process(array_obj_ref_333_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_333_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_333_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_rename
    process(LSHR_u64_u64_396_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_396_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_resize
    process(LSHR_u64_u64_396_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_396_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_root_address_inst
    process(array_obj_ref_397_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_397_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_397_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_addr_0
    process(ptr_deref_338_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_base_resize
    process(fetch_addr_335) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_335;
      ov := iv(13 downto 0);
      ptr_deref_338_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_gather_scatter
    process(ptr_deref_338_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_data_0;
      ov(63 downto 0) := iv;
      my_fetch_339 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_root_address_inst
    process(ptr_deref_338_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_addr_0
    process(ptr_deref_406_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_base_resize
    process(fetch_addr_399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_399;
      ov := iv(13 downto 0);
      ptr_deref_406_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_gather_scatter
    process(ptr_deref_406_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_data_0;
      ov(63 downto 0) := iv;
      fv_407 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_root_address_inst
    process(ptr_deref_406_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_350_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_425_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_350_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_350_branch_req_0,
          ack0 => do_while_stmt_350_branch_ack_0,
          ack1 => do_while_stmt_350_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_373_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_352, konst_372_wire_constant, tmp_var);
      nmycount_374 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_365_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_352, konst_364_wire_constant, tmp_var);
      AND_u64_u64_365_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_387_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_374, konst_386_wire_constant, tmp_var);
      AND_u64_u64_387_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_343_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_342_wire_constant, tmp_var);
      first_fill_344 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_389_inst
    process(AND_u64_u64_387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_387_wire, konst_388_wire_constant, tmp_var);
      fn_390 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_327_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_326_wire_constant, tmp_var);
      sh_start_328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_378_inst
    process(fetch_val_356, my_num1_369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_356, my_num1_369, tmp_var);
      LSHR_u64_u64_378_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_396_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_374, konst_395_wire_constant, tmp_var);
      LSHR_u64_u64_396_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_368_inst
    process(SUB_u64_u64_366_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_366_wire, konst_367_wire_constant, tmp_var);
      my_num1_369 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_366_inst
    process(konst_362_wire_constant, AND_u64_u64_365_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_362_wire_constant, AND_u64_u64_365_wire, tmp_var);
      SUB_u64_u64_366_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_424_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_423_wire_constant, tmp_var);
      SUB_u64_u64_424_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_431_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_431_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_425_inst
    process(mycount_352, SUB_u64_u64_424_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_352, SUB_u64_u64_424_wire, tmp_var);
      ULT_u64_u1_425_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_333_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_332_scaled;
      array_obj_ref_333_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_333_index_offset_req_0;
      array_obj_ref_333_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_333_index_offset_req_1;
      array_obj_ref_333_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_397_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_396_scaled;
      array_obj_ref_397_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_397_index_offset_req_0;
      array_obj_ref_397_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_397_index_offset_req_1;
      array_obj_ref_397_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_338_load_0 ptr_deref_406_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_338_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_406_load_0_req_0;
      ptr_deref_338_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_406_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_338_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_406_load_0_req_1;
      ptr_deref_338_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_406_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_388_delayed_7_0_402(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_338_word_address_0 & ptr_deref_406_word_address_0;
      ptr_deref_338_data_0 <= data_out(127 downto 64);
      ptr_deref_406_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_347_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_0;
      RPIPE_input_done_pipe_347_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_1;
      RPIPE_input_done_pipe_347_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_344(0);
      start_next_348 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_381_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_0;
      WPIPE_kernel_pipe1_381_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_1;
      WPIPE_kernel_pipe1_381_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val_380;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_size_pipe_428_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_0;
      WPIPE_size_pipe_428_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_1;
      WPIPE_size_pipe_428_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= first_fill_344(0);
      data_in <= type_cast_432_wire;
      size_pipe_write_1_gI: SplitGuardInterface generic map(name => "size_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_318_load_0_req_0 : boolean;
  signal LOAD_count_318_load_0_ack_0 : boolean;
  signal LOAD_count_318_load_0_req_1 : boolean;
  signal LOAD_count_318_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_319/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_sample_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_update_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/cr
      -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_1); -- 
    rr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_sample_completed_
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/ra
      -- 
    ra_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_0, ack => timer_CP_637_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_319/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_update_completed_
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_ack
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_1, ack => timer_CP_637_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_318_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_318_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_318_word_address_0 <= "0";
    -- equivalence LOAD_count_318_gather_scatter
    process(LOAD_count_318_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_318_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_318_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_318_load_0_req_0;
      LOAD_count_318_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_318_load_0_req_1;
      LOAD_count_318_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_318_word_address_0;
      LOAD_count_318_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_4576_start: Boolean;
  signal timerDaemon_CP_4576_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_2002_branch_req_0 : boolean;
  signal phi_stmt_2004_req_1 : boolean;
  signal phi_stmt_2004_req_0 : boolean;
  signal phi_stmt_2004_ack_0 : boolean;
  signal ADD_u64_u64_2010_inst_req_0 : boolean;
  signal ADD_u64_u64_2010_inst_ack_0 : boolean;
  signal ADD_u64_u64_2010_inst_req_1 : boolean;
  signal ADD_u64_u64_2010_inst_ack_1 : boolean;
  signal STORE_count_2012_store_0_req_0 : boolean;
  signal STORE_count_2012_store_0_ack_0 : boolean;
  signal STORE_count_2012_store_0_req_1 : boolean;
  signal STORE_count_2012_store_0_ack_1 : boolean;
  signal do_while_stmt_2002_branch_ack_0 : boolean;
  signal do_while_stmt_2002_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_4576_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4576_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_4576_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4576_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_4576: Block -- control-path 
    signal timerDaemon_CP_4576_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_4576_elements(0) <= timerDaemon_CP_4576_start;
    timerDaemon_CP_4576_symbol <= timerDaemon_CP_4576_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2001/$entry
      -- CP-element group 0: 	 branch_block_stmt_2001/branch_block_stmt_2001__entry__
      -- CP-element group 0: 	 branch_block_stmt_2001/do_while_stmt_2002__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2001/$exit
      -- CP-element group 1: 	 branch_block_stmt_2001/branch_block_stmt_2001__exit__
      -- CP-element group 1: 	 branch_block_stmt_2001/do_while_stmt_2002__exit__
      -- 
    timerDaemon_CP_4576_elements(1) <= timerDaemon_CP_4576_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2001/do_while_stmt_2002/$entry
      -- CP-element group 2: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002__entry__
      -- 
    timerDaemon_CP_4576_elements(2) <= timerDaemon_CP_4576_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002__exit__
      -- 
    -- Element group timerDaemon_CP_4576_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_back
      -- 
    -- Element group timerDaemon_CP_4576_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2001/do_while_stmt_2002/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_taken/$entry
      -- 
    timerDaemon_CP_4576_elements(5) <= timerDaemon_CP_4576_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_body_done
      -- 
    timerDaemon_CP_4576_elements(6) <= timerDaemon_CP_4576_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_4576_elements(7) <= timerDaemon_CP_4576_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_4576_elements(8) <= timerDaemon_CP_4576_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	31 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_4576_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/condition_evaluated
      -- 
    condition_evaluated_4600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(10), ack => do_while_stmt_2002_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(15) & timerDaemon_CP_4576_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(12) & timerDaemon_CP_4576_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(9) & timerDaemon_CP_4576_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(9) & timerDaemon_CP_4576_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_4576_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_4576_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_loopback_trigger
      -- 
    timerDaemon_CP_4576_elements(16) <= timerDaemon_CP_4576_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_loopback_sample_req_ps
      -- 
    phi_stmt_2004_loopback_sample_req_4615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2004_loopback_sample_req_4615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(17), ack => phi_stmt_2004_req_1); -- 
    -- Element group timerDaemon_CP_4576_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_entry_trigger
      -- 
    timerDaemon_CP_4576_elements(18) <= timerDaemon_CP_4576_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_entry_sample_req_ps
      -- 
    phi_stmt_2004_entry_sample_req_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2004_entry_sample_req_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(19), ack => phi_stmt_2004_req_0); -- 
    -- Element group timerDaemon_CP_4576_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/phi_stmt_2004_phi_mux_ack_ps
      -- 
    phi_stmt_2004_phi_mux_ack_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2004_ack_0, ack => timerDaemon_CP_4576_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_sample_completed_
      -- 
    -- Element group timerDaemon_CP_4576_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_update_start_
      -- 
    -- Element group timerDaemon_CP_4576_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_update_completed__ps
      -- 
    timerDaemon_CP_4576_elements(23) <= timerDaemon_CP_4576_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/type_cast_2007_update_completed_
      -- 
    -- Element group timerDaemon_CP_4576_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_4576_elements(22), ack => timerDaemon_CP_4576_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_4576_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_update_start__ps
      -- 
    -- Element group timerDaemon_CP_4576_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Sample/rr
      -- 
    rr_4642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(27), ack => ADD_u64_u64_2010_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(25) & timerDaemon_CP_4576_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Update/cr
      -- 
    cr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(28), ack => ADD_u64_u64_2010_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(26) & timerDaemon_CP_4576_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Sample/ra
      -- 
    ra_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2010_inst_ack_0, ack => timerDaemon_CP_4576_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/ADD_u64_u64_2010_Update/ca
      -- 
    ca_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2010_inst_ack_1, ack => timerDaemon_CP_4576_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/STORE_count_2012_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/STORE_count_2012_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/STORE_count_2012_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/STORE_count_2012_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/word_access_start/word_0/rr
      -- 
    rr_4670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(31), ack => STORE_count_2012_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(9) & timerDaemon_CP_4576_elements(15) & timerDaemon_CP_4576_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/word_access_complete/word_0/cr
      -- 
    cr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4576_elements(32), ack => STORE_count_2012_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_4576_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Sample/word_access_start/word_0/ra
      -- 
    ra_4671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2012_store_0_ack_0, ack => timerDaemon_CP_4576_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/STORE_count_2012_Update/word_access_complete/word_0/ca
      -- 
    ca_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2012_store_0_ack_1, ack => timerDaemon_CP_4576_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_4576_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_4576_elements(9), ack => timerDaemon_CP_4576_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_2001/do_while_stmt_2002/do_while_stmt_2002_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4576_elements(14) & timerDaemon_CP_4576_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4576_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_exit/ack
      -- 
    ack_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2002_branch_ack_0, ack => timerDaemon_CP_4576_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_2001/do_while_stmt_2002/loop_taken/ack
      -- 
    ack_4691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2002_branch_ack_1, ack => timerDaemon_CP_4576_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2001/do_while_stmt_2002/$exit
      -- 
    timerDaemon_CP_4576_elements(39) <= timerDaemon_CP_4576_elements(3);
    timerDaemon_do_while_stmt_2002_terminator_4692: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2002_terminator_4692", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_4576_elements(6),loop_continue => timerDaemon_CP_4576_elements(38),loop_terminate => timerDaemon_CP_4576_elements(37),loop_back => timerDaemon_CP_4576_elements(4),loop_exit => timerDaemon_CP_4576_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2004_phi_seq_4649_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_4576_elements(18);
      timerDaemon_CP_4576_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_4576_elements(21);
      timerDaemon_CP_4576_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_4576_elements(23);
      timerDaemon_CP_4576_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_4576_elements(16);
      timerDaemon_CP_4576_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_4576_elements(29);
      timerDaemon_CP_4576_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_4576_elements(30);
      timerDaemon_CP_4576_elements(17) <= phi_mux_reqs(1);
      phi_stmt_2004_phi_seq_4649 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_2004_phi_seq_4649") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_4576_elements(11), 
          phi_sample_ack => timerDaemon_CP_4576_elements(14), 
          phi_update_req => timerDaemon_CP_4576_elements(13), 
          phi_update_ack => timerDaemon_CP_4576_elements(15), 
          phi_mux_ack => timerDaemon_CP_4576_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4601_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_4576_elements(7);
        preds(1)  <= timerDaemon_CP_4576_elements(8);
        entry_tmerge_4601 : transition_merge -- 
          generic map(name => " entry_tmerge_4601")
          port map (preds => preds, symbol_out => timerDaemon_CP_4576_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_2010_wire : std_logic_vector(63 downto 0);
    signal STORE_count_2012_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_2012_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_2009_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2016_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_2004 : std_logic_vector(63 downto 0);
    signal type_cast_2007_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_2012_word_address_0 <= "0";
    konst_2009_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2016_wire_constant <= "1";
    type_cast_2007_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2004: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2007_wire_constant & ADD_u64_u64_2010_wire;
      req <= phi_stmt_2004_req_0 & phi_stmt_2004_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2004",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2004_ack_0,
          idata => idata,
          odata => ncount_2004,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2004
    -- equivalence STORE_count_2012_gather_scatter
    process(ncount_2004) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_2004;
      ov(63 downto 0) := iv;
      STORE_count_2012_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_2002_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2016_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2002_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2002_branch_req_0,
          ack0 => do_while_stmt_2002_branch_ack_0,
          ack1 => do_while_stmt_2002_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_2010_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_2004;
      ADD_u64_u64_2010_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2010_inst_req_0;
      ADD_u64_u64_2010_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2010_inst_req_1;
      ADD_u64_u64_2010_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_2012_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_2012_store_0_req_0;
      STORE_count_2012_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_2012_store_0_req_1;
      STORE_count_2012_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_2012_word_address_0;
      data_in <= STORE_count_2012_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(127 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(127 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(127 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(127 downto 64);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(63 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 128,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
