-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_59_branch_req_0 : boolean;
  signal if_stmt_59_branch_ack_1 : boolean;
  signal if_stmt_59_branch_ack_0 : boolean;
  signal type_cast_68_inst_req_0 : boolean;
  signal type_cast_68_inst_ack_0 : boolean;
  signal type_cast_68_inst_req_1 : boolean;
  signal type_cast_68_inst_ack_1 : boolean;
  signal array_obj_ref_84_index_offset_req_0 : boolean;
  signal array_obj_ref_84_index_offset_ack_0 : boolean;
  signal array_obj_ref_84_index_offset_req_1 : boolean;
  signal array_obj_ref_84_index_offset_ack_1 : boolean;
  signal addr_of_85_final_reg_req_0 : boolean;
  signal addr_of_85_final_reg_ack_0 : boolean;
  signal addr_of_85_final_reg_req_1 : boolean;
  signal addr_of_85_final_reg_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_177_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_177_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_177_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_177_inst_ack_1 : boolean;
  signal ptr_deref_89_load_0_req_0 : boolean;
  signal ptr_deref_89_load_0_ack_0 : boolean;
  signal ptr_deref_89_load_0_req_1 : boolean;
  signal ptr_deref_89_load_0_ack_1 : boolean;
  signal type_cast_93_inst_req_0 : boolean;
  signal type_cast_93_inst_ack_0 : boolean;
  signal type_cast_93_inst_req_1 : boolean;
  signal type_cast_93_inst_ack_1 : boolean;
  signal type_cast_103_inst_req_0 : boolean;
  signal type_cast_103_inst_ack_0 : boolean;
  signal type_cast_103_inst_req_1 : boolean;
  signal type_cast_103_inst_ack_1 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal type_cast_123_inst_req_0 : boolean;
  signal type_cast_123_inst_ack_0 : boolean;
  signal type_cast_123_inst_req_1 : boolean;
  signal type_cast_123_inst_ack_1 : boolean;
  signal type_cast_133_inst_req_0 : boolean;
  signal type_cast_133_inst_ack_0 : boolean;
  signal type_cast_133_inst_req_1 : boolean;
  signal type_cast_133_inst_ack_1 : boolean;
  signal type_cast_143_inst_req_0 : boolean;
  signal type_cast_143_inst_ack_0 : boolean;
  signal type_cast_143_inst_req_1 : boolean;
  signal type_cast_143_inst_ack_1 : boolean;
  signal type_cast_153_inst_req_0 : boolean;
  signal type_cast_153_inst_ack_0 : boolean;
  signal type_cast_153_inst_req_1 : boolean;
  signal type_cast_153_inst_ack_1 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_174_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_174_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_174_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_174_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_180_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_180_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_180_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_180_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_183_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_183_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_183_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_183_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_186_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_186_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_186_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_186_inst_ack_1 : boolean;
  signal if_stmt_200_branch_req_0 : boolean;
  signal if_stmt_200_branch_ack_1 : boolean;
  signal if_stmt_200_branch_ack_0 : boolean;
  signal phi_stmt_72_req_0 : boolean;
  signal type_cast_78_inst_req_0 : boolean;
  signal type_cast_78_inst_ack_0 : boolean;
  signal type_cast_78_inst_req_1 : boolean;
  signal type_cast_78_inst_ack_1 : boolean;
  signal phi_stmt_72_req_1 : boolean;
  signal phi_stmt_72_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_39/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/branch_block_stmt_39__entry__
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_49_to_assign_stmt_58__entry__
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_49_to_assign_stmt_58__exit__
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59__entry__
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_49_to_assign_stmt_58/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/assign_stmt_49_to_assign_stmt_58/$exit
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_39/R_cmp68_60_place
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_39/if_stmt_59_else_link/$entry
      -- 
    branch_req_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => if_stmt_59_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_39/merge_stmt_65__exit__
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69__entry__
      -- CP-element group 1: 	 branch_block_stmt_39/if_stmt_59_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_39/if_stmt_59_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_39/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/$entry
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_update_start_
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_39/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_39/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_39/merge_stmt_65_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_39/merge_stmt_65_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_39/merge_stmt_65_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_39/merge_stmt_65_PhiAck/dummy
      -- 
    if_choice_transition_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_59_branch_ack_1, ack => sendOutput_CP_26_elements(1)); -- 
    rr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_68_inst_req_0); -- 
    cr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_68_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_39/if_stmt_59_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_39/if_stmt_59_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_39/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_39/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_39/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_59_branch_ack_0, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Sample/ra
      -- 
    ra_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_69__exit__
      -- CP-element group 4: 	 branch_block_stmt_39/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_69/$exit
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_39/assign_stmt_69/type_cast_68_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/phi_stmt_72/$entry
      -- CP-element group 4: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/$entry
      -- 
    ca_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Sample/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_84_index_offset_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_request/req
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_84_index_offset_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(6), ack => addr_of_85_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_request/ack
      -- 
    ack_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_85_final_reg_ack_0, ack => sendOutput_CP_26_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/word_access_start/word_0/rr
      -- 
    ack_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_85_final_reg_ack_1, ack => sendOutput_CP_26_elements(8)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(8), ack => ptr_deref_89_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Sample/word_access_start/word_0/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_89_load_0_ack_0, ack => sendOutput_CP_26_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/ptr_deref_89_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/ptr_deref_89_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/ptr_deref_89_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/ptr_deref_89_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_89_load_0_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_123_inst_req_0); -- 
    rr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_133_inst_req_0); -- 
    rr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_143_inst_req_0); -- 
    rr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_153_inst_req_0); -- 
    rr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_163_inst_req_0); -- 
    rr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_93_inst_req_0); -- 
    rr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_113_inst_req_0); -- 
    rr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_103_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Sample/ra
      -- 
    ra_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Update/ca
      -- 
    ca_205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_1, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Sample/ra
      -- 
    ra_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_103_inst_ack_0, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Update/ca
      -- 
    ca_219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_103_inst_ack_1, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Sample/ra
      -- 
    ra_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => sendOutput_CP_26_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Update/ca
      -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Sample/ra
      -- 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_123_inst_ack_0, ack => sendOutput_CP_26_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Update/ca
      -- 
    ca_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_123_inst_ack_1, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Sample/ra
      -- 
    ra_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_133_inst_ack_0, ack => sendOutput_CP_26_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Update/ca
      -- 
    ca_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_133_inst_ack_1, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Sample/ra
      -- 
    ra_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_0, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Update/ca
      -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_1, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Sample/ra
      -- 
    ra_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_0, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Update/ca
      -- 
    ca_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_1, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Sample/ra
      -- 
    ra_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Sample/req
      -- 
    ca_303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => sendOutput_CP_26_elements(26)); -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(26), ack => WPIPE_zeropad_output_pipe_165_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_update_start_
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Update/req
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_165_inst_ack_0, ack => sendOutput_CP_26_elements(27)); -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(27), ack => WPIPE_zeropad_output_pipe_165_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_165_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_165_inst_ack_1, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Sample/req
      -- 
    req_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(29), ack => WPIPE_zeropad_output_pipe_168_inst_req_0); -- 
    sendOutput_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(24) & sendOutput_CP_26_elements(28);
      gj_sendOutput_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_update_start_
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Update/req
      -- 
    ack_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_168_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(30), ack => WPIPE_zeropad_output_pipe_168_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_168_Update/ack
      -- 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_168_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	22 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Sample/req
      -- 
    req_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(32), ack => WPIPE_zeropad_output_pipe_171_inst_req_0); -- 
    sendOutput_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(22) & sendOutput_CP_26_elements(31);
      gj_sendOutput_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_update_start_
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Update/req
      -- 
    ack_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_171_inst_ack_0, ack => sendOutput_CP_26_elements(33)); -- 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(33), ack => WPIPE_zeropad_output_pipe_171_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_171_Update/ack
      -- 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_171_inst_ack_1, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	20 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Sample/req
      -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_174_inst_req_0); -- 
    sendOutput_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(20) & sendOutput_CP_26_elements(34);
      gj_sendOutput_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_update_start_
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Update/req
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_174_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_174_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_174_Update/ack
      -- 
    ack_359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_174_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_sample_start_
      -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_177_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(18) & sendOutput_CP_26_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_update_start_
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Update/req
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_177_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_177_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_177_Update/ack
      -- 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_177_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Sample/req
      -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_180_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(16) & sendOutput_CP_26_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_update_start_
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Update/req
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_180_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_180_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_180_Update/ack
      -- 
    ack_387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_180_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	14 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Sample/req
      -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_183_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(43) & sendOutput_CP_26_elements(14);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_update_start_
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Update/req
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_183_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_183_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_183_Update/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_183_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	12 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_186_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(12) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_update_start_
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Update/req
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_186_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_186_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/WPIPE_zeropad_output_pipe_186_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_186_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199__exit__
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200__entry__
      -- CP-element group 50: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/$exit
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_39/R_exitcond2_201_place
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_39/if_stmt_200_else_link/$entry
      -- 
    branch_req_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => if_stmt_200_branch_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(5) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_39/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_39/merge_stmt_206__exit__
      -- CP-element group 51: 	 branch_block_stmt_39/if_stmt_200_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_39/if_stmt_200_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_39/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_39/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_39/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_39/merge_stmt_206_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_39/merge_stmt_206_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_39/merge_stmt_206_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_39/merge_stmt_206_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_39/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_39/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_200_branch_ack_1, ack => sendOutput_CP_26_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_39/if_stmt_200_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_39/if_stmt_200_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Update/cr
      -- 
    else_choice_transition_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_200_branch_ack_0, ack => sendOutput_CP_26_elements(52)); -- 
    rr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_78_inst_req_0); -- 
    cr_481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_78_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/phi_stmt_72/$exit
      -- CP-element group 53: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_76_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_39/bbx_xnph_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_req
      -- 
    phi_stmt_72_req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_72_req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => phi_stmt_72_req_0); -- 
    -- Element group sendOutput_CP_26_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(4), ack => sendOutput_CP_26_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Sample/ra
      -- 
    ra_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_78_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/Update/ca
      -- 
    ca_482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_78_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/$exit
      -- CP-element group 56: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/$exit
      -- CP-element group 56: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_sources/type_cast_78/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_39/forx_xbody_forx_xbody_PhiReq/phi_stmt_72/phi_stmt_72_req
      -- 
    phi_stmt_72_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_72_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => phi_stmt_72_req_1); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(54) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_39/merge_stmt_71_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_39/merge_stmt_71_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(57) <= OrReduce(sendOutput_CP_26_elements(53) & sendOutput_CP_26_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	24 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_39/merge_stmt_71__exit__
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199__entry__
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/array_obj_ref_84_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/addr_of_85_complete/req
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/ptr_deref_89_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_93_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_103_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_113_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_123_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_133_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_143_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_153_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_update_start_
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_39/assign_stmt_86_to_assign_stmt_199/type_cast_163_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_39/merge_stmt_71_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_39/merge_stmt_71_PhiAck/phi_stmt_72_ack
      -- 
    phi_stmt_72_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_72_ack_0, ack => sendOutput_CP_26_elements(58)); -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_84_index_offset_req_0); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_84_index_offset_req_1); -- 
    req_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => addr_of_85_final_reg_req_1); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => ptr_deref_89_load_0_req_1); -- 
    cr_204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_93_inst_req_1); -- 
    cr_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_103_inst_req_1); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_113_inst_req_1); -- 
    cr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_123_inst_req_1); -- 
    cr_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_133_inst_req_1); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_143_inst_req_1); -- 
    cr_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_153_inst_req_1); -- 
    cr_302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_163_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_208__exit__
      -- CP-element group 59: 	 branch_block_stmt_39/return__
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_210__exit__
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_39/$exit
      -- CP-element group 59: 	 branch_block_stmt_39/branch_block_stmt_39__exit__
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_208_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_208_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_208_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_208_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_39/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_39/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_210_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_210_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_210_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_39/merge_stmt_210_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(59) <= OrReduce(sendOutput_CP_26_elements(2) & sendOutput_CP_26_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_47_wire : std_logic_vector(31 downto 0);
    signal R_indvar_83_resized : std_logic_vector(13 downto 0);
    signal R_indvar_83_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_84_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_84_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_84_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_84_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_84_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_84_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_86 : std_logic_vector(31 downto 0);
    signal cmp68_58 : std_logic_vector(0 downto 0);
    signal conv12_104 : std_logic_vector(7 downto 0);
    signal conv18_114 : std_logic_vector(7 downto 0);
    signal conv24_124 : std_logic_vector(7 downto 0);
    signal conv30_134 : std_logic_vector(7 downto 0);
    signal conv36_144 : std_logic_vector(7 downto 0);
    signal conv42_154 : std_logic_vector(7 downto 0);
    signal conv48_164 : std_logic_vector(7 downto 0);
    signal conv_94 : std_logic_vector(7 downto 0);
    signal exitcond2_199 : std_logic_vector(0 downto 0);
    signal indvar_72 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_194 : std_logic_vector(63 downto 0);
    signal ptr_deref_89_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_89_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_89_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_89_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_89_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_110 : std_logic_vector(63 downto 0);
    signal shr21_120 : std_logic_vector(63 downto 0);
    signal shr27_130 : std_logic_vector(63 downto 0);
    signal shr33_140 : std_logic_vector(63 downto 0);
    signal shr39_150 : std_logic_vector(63 downto 0);
    signal shr45_160 : std_logic_vector(63 downto 0);
    signal shr67_49 : std_logic_vector(31 downto 0);
    signal shr9_100 : std_logic_vector(63 downto 0);
    signal tmp1_69 : std_logic_vector(63 downto 0);
    signal tmp4_90 : std_logic_vector(63 downto 0);
    signal type_cast_108_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_138_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_148_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_158_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_192_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_43_wire : std_logic_vector(31 downto 0);
    signal type_cast_46_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_52_wire : std_logic_vector(31 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_76_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_78_wire : std_logic_vector(63 downto 0);
    signal type_cast_98_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_84_constant_part_of_offset <= "00000000000000";
    array_obj_ref_84_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_84_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_84_resized_base_address <= "00000000000000";
    ptr_deref_89_word_offset_0 <= "00000000000000";
    type_cast_108_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_118_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_128_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_138_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_148_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_158_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_192_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_46_wire_constant <= "00000000000000000000000000000010";
    type_cast_55_wire_constant <= "00000000000000000000000000000000";
    type_cast_76_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_98_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    phi_stmt_72: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_76_wire_constant & type_cast_78_wire;
      req <= phi_stmt_72_req_0 & phi_stmt_72_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_72",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_72_ack_0,
          idata => idata,
          odata => indvar_72,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_72
    addr_of_85_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_85_final_reg_req_0;
      addr_of_85_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_85_final_reg_req_1;
      addr_of_85_final_reg_ack_1<= rack(0);
      addr_of_85_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_85_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_84_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_86,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_103_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_103_inst_req_0;
      type_cast_103_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_103_inst_req_1;
      type_cast_103_inst_ack_1<= rack(0);
      type_cast_103_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_103_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_123_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_123_inst_req_0;
      type_cast_123_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_123_inst_req_1;
      type_cast_123_inst_ack_1<= rack(0);
      type_cast_123_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_123_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_133_inst_req_0;
      type_cast_133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_133_inst_req_1;
      type_cast_133_inst_ack_1<= rack(0);
      type_cast_133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_133_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_143_inst_req_0;
      type_cast_143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_143_inst_req_1;
      type_cast_143_inst_ack_1<= rack(0);
      type_cast_143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_153_inst_req_0;
      type_cast_153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_153_inst_req_1;
      type_cast_153_inst_ack_1<= rack(0);
      type_cast_153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_150,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_154,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_43_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := size_buffer(31 downto 0);
      type_cast_43_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_48_inst
    process(ASHR_i32_i32_47_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_47_wire(31 downto 0);
      shr67_49 <= tmp_var; -- 
    end process;
    -- interlock type_cast_52_inst
    process(shr67_49) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := shr67_49(31 downto 0);
      type_cast_52_wire <= tmp_var; -- 
    end process;
    type_cast_68_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_68_inst_req_0;
      type_cast_68_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_68_inst_req_1;
      type_cast_68_inst_ack_1<= rack(0);
      type_cast_68_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_68_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr67_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_69,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_78_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_78_inst_req_0;
      type_cast_78_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_78_inst_req_1;
      type_cast_78_inst_ack_1<= rack(0);
      type_cast_78_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_78_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_78_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_93_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_93_inst_req_0;
      type_cast_93_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_93_inst_req_1;
      type_cast_93_inst_ack_1<= rack(0);
      type_cast_93_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_93_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_90,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_94,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_84_index_1_rename
    process(R_indvar_83_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_83_resized;
      ov(13 downto 0) := iv;
      R_indvar_83_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_84_index_1_resize
    process(indvar_72) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_72;
      ov := iv(13 downto 0);
      R_indvar_83_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_84_root_address_inst
    process(array_obj_ref_84_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_84_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_84_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_89_addr_0
    process(ptr_deref_89_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_89_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_89_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_89_base_resize
    process(arrayidx_86) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_86;
      ov := iv(13 downto 0);
      ptr_deref_89_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_89_gather_scatter
    process(ptr_deref_89_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_89_data_0;
      ov(63 downto 0) := iv;
      tmp4_90 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_89_root_address_inst
    process(ptr_deref_89_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_89_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_89_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_200_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_199;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_200_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_200_branch_req_0,
          ack0 => if_stmt_200_branch_ack_0,
          ack1 => if_stmt_200_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_59_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_58;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_59_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_59_branch_req_0,
          ack0 => if_stmt_59_branch_ack_0,
          ack1 => if_stmt_59_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_193_inst
    process(indvar_72) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_72, type_cast_192_wire_constant, tmp_var);
      indvarx_xnext_194 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_47_inst
    process(type_cast_43_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_43_wire, type_cast_46_wire_constant, tmp_var);
      ASHR_i32_i32_47_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_198_inst
    process(indvarx_xnext_194, tmp1_69) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_194, tmp1_69, tmp_var);
      exitcond2_199 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_109_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_108_wire_constant, tmp_var);
      shr15_110 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_119_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_118_wire_constant, tmp_var);
      shr21_120 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_129_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_128_wire_constant, tmp_var);
      shr27_130 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_139_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_138_wire_constant, tmp_var);
      shr33_140 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_149_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_148_wire_constant, tmp_var);
      shr39_150 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_159_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_158_wire_constant, tmp_var);
      shr45_160 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_99_inst
    process(tmp4_90) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_90, type_cast_98_wire_constant, tmp_var);
      shr9_100 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_56_inst
    process(type_cast_52_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_52_wire, type_cast_55_wire_constant, tmp_var);
      cmp68_58 <= tmp_var; --
    end process;
    -- shared split operator group (11) : array_obj_ref_84_index_offset 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_83_scaled;
      array_obj_ref_84_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_84_index_offset_req_0;
      array_obj_ref_84_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_84_index_offset_req_1;
      array_obj_ref_84_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared load operator group (0) : ptr_deref_89_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_89_load_0_req_0;
      ptr_deref_89_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_89_load_0_req_1;
      ptr_deref_89_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_89_word_address_0;
      ptr_deref_89_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_165_inst WPIPE_zeropad_output_pipe_168_inst WPIPE_zeropad_output_pipe_171_inst WPIPE_zeropad_output_pipe_174_inst WPIPE_zeropad_output_pipe_177_inst WPIPE_zeropad_output_pipe_180_inst WPIPE_zeropad_output_pipe_183_inst WPIPE_zeropad_output_pipe_186_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_165_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_168_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_171_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_174_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_177_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_180_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_183_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_186_inst_req_0;
      WPIPE_zeropad_output_pipe_165_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_168_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_171_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_174_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_177_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_180_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_183_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_186_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_165_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_168_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_171_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_174_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_177_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_180_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_183_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_186_inst_req_1;
      WPIPE_zeropad_output_pipe_165_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_168_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_171_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_174_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_177_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_180_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_183_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_186_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv48_164 & conv42_154 & conv36_144 & conv30_134 & conv24_124 & conv18_114 & conv12_104 & conv_94;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_520_start: Boolean;
  signal timer_CP_520_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_216_load_0_ack_1 : boolean;
  signal LOAD_count_216_load_0_req_1 : boolean;
  signal LOAD_count_216_load_0_ack_0 : boolean;
  signal LOAD_count_216_load_0_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_520_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_520: Block -- control-path 
    signal timer_CP_520_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_520_elements(0) <= timer_CP_520_start;
    timer_CP_520_symbol <= timer_CP_520_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_update_start_
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_sample_start_
      -- CP-element group 0: 	 assign_stmt_217/$entry
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Update/$entry
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_217/LOAD_count_216_Sample/word_access_start/$entry
      -- CP-element group 0: 	 $entry
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_216_load_0_req_1); -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_216_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_217/LOAD_count_216_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_217/LOAD_count_216_sample_completed_
      -- CP-element group 1: 	 assign_stmt_217/LOAD_count_216_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_217/LOAD_count_216_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_217/LOAD_count_216_Sample/word_access_start/$exit
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_216_load_0_ack_0, ack => timer_CP_520_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/LOAD_count_216_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/LOAD_count_216_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_217/$exit
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_update_completed_
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/$exit
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/LOAD_count_216_Merge/merge_ack
      -- CP-element group 2: 	 assign_stmt_217/LOAD_count_216_Update/LOAD_count_216_Merge/merge_req
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_216_load_0_ack_1, ack => timer_CP_520_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_216_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_216_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_216_word_address_0 <= "0";
    -- equivalence LOAD_count_216_gather_scatter
    process(LOAD_count_216_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_216_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_216_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_216_load_0_req_0;
      LOAD_count_216_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_216_load_0_req_1;
      LOAD_count_216_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_216_word_address_0;
      LOAD_count_216_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block3_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block4_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block4_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block4_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block5_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block5_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block5_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block6_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block6_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block6_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block7_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block7_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block7_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block3_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block7_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block7_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block7_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    Block4_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block4_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block4_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block5_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block5_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block5_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block6_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block6_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block6_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_data : out  std_logic_vector(31 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_676_start: Boolean;
  signal zeropad3D_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_zeropad_input_pipe_250_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_253_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_598_inst_req_1 : boolean;
  signal WPIPE_Block4_starting_634_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_622_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_595_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_577_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_244_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_640_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_595_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_244_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_577_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_634_inst_req_1 : boolean;
  signal WPIPE_Block4_starting_619_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_571_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_559_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_562_inst_req_1 : boolean;
  signal WPIPE_Block5_starting_640_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_577_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_571_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_577_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_571_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_559_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_619_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_601_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_613_inst_req_0 : boolean;
  signal WPIPE_Block5_starting_640_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_241_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_259_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_241_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_259_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_595_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_574_inst_req_0 : boolean;
  signal WPIPE_Block5_starting_640_inst_req_1 : boolean;
  signal WPIPE_Block5_starting_646_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_595_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_592_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_634_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_592_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_628_inst_ack_1 : boolean;
  signal type_cast_273_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_568_inst_req_1 : boolean;
  signal type_cast_310_inst_ack_1 : boolean;
  signal type_cast_310_inst_req_0 : boolean;
  signal type_cast_310_inst_ack_0 : boolean;
  signal type_cast_310_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_601_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_247_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_646_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_247_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_592_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_604_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_601_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_601_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_247_inst_ack_0 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_ack_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal WPIPE_Block5_starting_649_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_265_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_265_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_req_1 : boolean;
  signal WPIPE_Block4_starting_625_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_250_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_562_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_256_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_256_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_256_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_256_inst_req_0 : boolean;
  signal type_cast_273_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_265_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_589_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_556_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_247_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_604_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_622_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_265_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_589_inst_req_1 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_259_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_259_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_556_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_253_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_241_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_634_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_253_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_241_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_562_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_562_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_262_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_628_inst_ack_0 : boolean;
  signal type_cast_314_inst_req_0 : boolean;
  signal type_cast_314_inst_ack_0 : boolean;
  signal type_cast_314_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_610_inst_ack_1 : boolean;
  signal type_cast_314_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_244_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_628_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_589_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_568_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_571_inst_req_0 : boolean;
  signal type_cast_277_inst_ack_1 : boolean;
  signal type_cast_277_inst_req_1 : boolean;
  signal type_cast_277_inst_req_0 : boolean;
  signal type_cast_277_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_625_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_244_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_592_inst_req_0 : boolean;
  signal if_stmt_301_branch_req_0 : boolean;
  signal WPIPE_Block2_starting_589_inst_req_0 : boolean;
  signal if_stmt_301_branch_ack_0 : boolean;
  signal if_stmt_301_branch_ack_1 : boolean;
  signal WPIPE_Block3_starting_598_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_253_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_628_inst_req_0 : boolean;
  signal type_cast_323_inst_req_0 : boolean;
  signal type_cast_323_inst_ack_0 : boolean;
  signal type_cast_323_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_610_inst_req_1 : boolean;
  signal type_cast_323_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_655_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_622_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_616_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_616_inst_req_1 : boolean;
  signal WPIPE_Block5_starting_649_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_586_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_646_inst_ack_0 : boolean;
  signal array_obj_ref_363_index_offset_req_0 : boolean;
  signal array_obj_ref_363_index_offset_ack_0 : boolean;
  signal array_obj_ref_363_index_offset_req_1 : boolean;
  signal array_obj_ref_363_index_offset_ack_1 : boolean;
  signal WPIPE_Block2_starting_586_inst_req_1 : boolean;
  signal WPIPE_Block5_starting_646_inst_req_0 : boolean;
  signal addr_of_364_final_reg_req_0 : boolean;
  signal WPIPE_Block3_starting_610_inst_ack_0 : boolean;
  signal addr_of_364_final_reg_ack_0 : boolean;
  signal addr_of_364_final_reg_req_1 : boolean;
  signal addr_of_364_final_reg_ack_1 : boolean;
  signal WPIPE_Block5_starting_655_inst_req_1 : boolean;
  signal WPIPE_Block4_starting_622_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_610_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_568_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_1 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_574_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_380_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_380_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_568_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_380_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_380_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_652_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_586_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_616_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_586_inst_req_0 : boolean;
  signal type_cast_384_inst_req_0 : boolean;
  signal type_cast_384_inst_ack_0 : boolean;
  signal type_cast_384_inst_req_1 : boolean;
  signal type_cast_384_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_398_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_398_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_398_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_398_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_652_inst_req_1 : boolean;
  signal WPIPE_Block4_starting_616_inst_req_0 : boolean;
  signal type_cast_402_inst_req_0 : boolean;
  signal type_cast_402_inst_ack_0 : boolean;
  signal type_cast_402_inst_req_1 : boolean;
  signal type_cast_402_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_637_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_655_inst_ack_0 : boolean;
  signal WPIPE_Block5_starting_637_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_416_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_416_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_416_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_416_inst_ack_1 : boolean;
  signal type_cast_420_inst_req_0 : boolean;
  signal type_cast_420_inst_ack_0 : boolean;
  signal type_cast_420_inst_req_1 : boolean;
  signal type_cast_420_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_655_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_434_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_434_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_434_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_434_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_631_inst_ack_1 : boolean;
  signal type_cast_438_inst_req_0 : boolean;
  signal type_cast_438_inst_ack_0 : boolean;
  signal type_cast_438_inst_req_1 : boolean;
  signal type_cast_438_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_637_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_452_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_452_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_452_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_452_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_631_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_583_inst_ack_1 : boolean;
  signal type_cast_456_inst_req_0 : boolean;
  signal type_cast_456_inst_ack_0 : boolean;
  signal type_cast_456_inst_req_1 : boolean;
  signal type_cast_456_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_649_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_637_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_470_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_607_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_470_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_470_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_470_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_652_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_631_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_583_inst_req_1 : boolean;
  signal type_cast_474_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_607_inst_req_1 : boolean;
  signal type_cast_474_inst_ack_0 : boolean;
  signal type_cast_474_inst_req_1 : boolean;
  signal type_cast_474_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_649_inst_req_1 : boolean;
  signal WPIPE_Block4_starting_619_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_488_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_488_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_488_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_488_inst_ack_1 : boolean;
  signal WPIPE_Block5_starting_652_inst_req_0 : boolean;
  signal WPIPE_Block4_starting_631_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_583_inst_ack_0 : boolean;
  signal type_cast_492_inst_req_0 : boolean;
  signal type_cast_492_inst_ack_0 : boolean;
  signal type_cast_492_inst_req_1 : boolean;
  signal type_cast_492_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_613_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_613_inst_req_1 : boolean;
  signal WPIPE_Block5_starting_643_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_607_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_583_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_598_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_574_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_607_inst_req_0 : boolean;
  signal WPIPE_Block5_starting_643_inst_req_1 : boolean;
  signal ptr_deref_500_store_0_req_0 : boolean;
  signal ptr_deref_500_store_0_ack_0 : boolean;
  signal WPIPE_Block3_starting_598_inst_req_0 : boolean;
  signal ptr_deref_500_store_0_req_1 : boolean;
  signal ptr_deref_500_store_0_ack_1 : boolean;
  signal WPIPE_Block2_starting_580_inst_ack_1 : boolean;
  signal WPIPE_Block4_starting_625_inst_ack_1 : boolean;
  signal if_stmt_514_branch_req_0 : boolean;
  signal WPIPE_Block2_starting_580_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_559_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_559_inst_req_1 : boolean;
  signal if_stmt_514_branch_ack_1 : boolean;
  signal if_stmt_514_branch_ack_0 : boolean;
  signal WPIPE_Block4_starting_619_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_574_inst_ack_0 : boolean;
  signal WPIPE_Block4_starting_625_inst_req_1 : boolean;
  signal call_stmt_525_call_req_0 : boolean;
  signal call_stmt_525_call_ack_0 : boolean;
  signal call_stmt_525_call_req_1 : boolean;
  signal call_stmt_525_call_ack_1 : boolean;
  signal WPIPE_Block1_starting_565_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_565_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_580_inst_ack_0 : boolean;
  signal type_cast_530_inst_req_0 : boolean;
  signal type_cast_530_inst_ack_0 : boolean;
  signal type_cast_530_inst_req_1 : boolean;
  signal type_cast_530_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_613_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_580_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_532_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_532_inst_ack_0 : boolean;
  signal WPIPE_Block5_starting_643_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_532_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_604_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_532_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_565_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_535_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_604_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_535_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_565_inst_req_0 : boolean;
  signal WPIPE_Block5_starting_643_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_535_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_535_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_538_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_538_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_538_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_538_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_541_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_541_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_541_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_541_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_544_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_544_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_544_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_544_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_547_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_547_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_547_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_547_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_550_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_550_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_550_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_550_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_553_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_553_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_553_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_553_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_556_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_556_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_658_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_658_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_658_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_658_inst_ack_1 : boolean;
  signal WPIPE_Block6_starting_661_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_661_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_661_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_661_inst_ack_1 : boolean;
  signal WPIPE_Block6_starting_664_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_664_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_664_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_664_inst_ack_1 : boolean;
  signal WPIPE_Block6_starting_667_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_667_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_667_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_667_inst_ack_1 : boolean;
  signal WPIPE_Block6_starting_670_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_670_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_670_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_670_inst_ack_1 : boolean;
  signal WPIPE_Block6_starting_673_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_673_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_673_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_673_inst_ack_1 : boolean;
  signal WPIPE_Block6_starting_676_inst_req_0 : boolean;
  signal WPIPE_Block6_starting_676_inst_ack_0 : boolean;
  signal WPIPE_Block6_starting_676_inst_req_1 : boolean;
  signal WPIPE_Block6_starting_676_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_679_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_679_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_679_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_679_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_682_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_682_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_682_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_682_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_685_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_685_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_685_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_685_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_688_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_688_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_688_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_688_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_691_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_691_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_691_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_691_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_694_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_694_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_694_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_694_inst_ack_1 : boolean;
  signal WPIPE_Block7_starting_697_inst_req_0 : boolean;
  signal WPIPE_Block7_starting_697_inst_ack_0 : boolean;
  signal WPIPE_Block7_starting_697_inst_req_1 : boolean;
  signal WPIPE_Block7_starting_697_inst_ack_1 : boolean;
  signal RPIPE_Block0_complete_702_inst_req_0 : boolean;
  signal RPIPE_Block0_complete_702_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_702_inst_req_1 : boolean;
  signal RPIPE_Block0_complete_702_inst_ack_1 : boolean;
  signal RPIPE_Block1_complete_705_inst_req_0 : boolean;
  signal RPIPE_Block1_complete_705_inst_ack_0 : boolean;
  signal RPIPE_Block1_complete_705_inst_req_1 : boolean;
  signal RPIPE_Block1_complete_705_inst_ack_1 : boolean;
  signal RPIPE_Block2_complete_708_inst_req_0 : boolean;
  signal RPIPE_Block2_complete_708_inst_ack_0 : boolean;
  signal RPIPE_Block2_complete_708_inst_req_1 : boolean;
  signal RPIPE_Block2_complete_708_inst_ack_1 : boolean;
  signal RPIPE_Block3_complete_711_inst_req_0 : boolean;
  signal RPIPE_Block3_complete_711_inst_ack_0 : boolean;
  signal RPIPE_Block3_complete_711_inst_req_1 : boolean;
  signal RPIPE_Block3_complete_711_inst_ack_1 : boolean;
  signal RPIPE_Block4_complete_714_inst_req_0 : boolean;
  signal RPIPE_Block4_complete_714_inst_ack_0 : boolean;
  signal RPIPE_Block4_complete_714_inst_req_1 : boolean;
  signal RPIPE_Block4_complete_714_inst_ack_1 : boolean;
  signal RPIPE_Block5_complete_717_inst_req_0 : boolean;
  signal RPIPE_Block5_complete_717_inst_ack_0 : boolean;
  signal RPIPE_Block5_complete_717_inst_req_1 : boolean;
  signal RPIPE_Block5_complete_717_inst_ack_1 : boolean;
  signal RPIPE_Block6_complete_720_inst_req_0 : boolean;
  signal RPIPE_Block6_complete_720_inst_ack_0 : boolean;
  signal RPIPE_Block6_complete_720_inst_req_1 : boolean;
  signal RPIPE_Block6_complete_720_inst_ack_1 : boolean;
  signal RPIPE_Block7_complete_723_inst_req_0 : boolean;
  signal RPIPE_Block7_complete_723_inst_ack_0 : boolean;
  signal RPIPE_Block7_complete_723_inst_req_1 : boolean;
  signal RPIPE_Block7_complete_723_inst_ack_1 : boolean;
  signal call_stmt_727_call_req_0 : boolean;
  signal call_stmt_727_call_ack_0 : boolean;
  signal call_stmt_727_call_req_1 : boolean;
  signal call_stmt_727_call_ack_1 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_738_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_738_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_738_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_738_inst_ack_1 : boolean;
  signal type_cast_744_inst_req_0 : boolean;
  signal type_cast_744_inst_ack_0 : boolean;
  signal type_cast_744_inst_req_1 : boolean;
  signal type_cast_744_inst_ack_1 : boolean;
  signal type_cast_748_inst_req_0 : boolean;
  signal type_cast_748_inst_ack_0 : boolean;
  signal type_cast_748_inst_req_1 : boolean;
  signal type_cast_748_inst_ack_1 : boolean;
  signal type_cast_752_inst_req_0 : boolean;
  signal type_cast_752_inst_ack_0 : boolean;
  signal type_cast_752_inst_req_1 : boolean;
  signal type_cast_752_inst_ack_1 : boolean;
  signal call_stmt_765_call_req_0 : boolean;
  signal call_stmt_765_call_ack_0 : boolean;
  signal call_stmt_765_call_req_1 : boolean;
  signal call_stmt_765_call_ack_1 : boolean;
  signal phi_stmt_351_req_0 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal phi_stmt_351_req_1 : boolean;
  signal phi_stmt_351_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_676: Block -- control-path 
    signal zeropad3D_CP_676_elements: BooleanArray(232 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_676_elements(0) <= zeropad3D_CP_676_start;
    zeropad3D_CP_676_symbol <= zeropad3D_CP_676_elements(225);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	22 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300__entry__
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/$entry
      -- CP-element group 0: 	 branch_block_stmt_239/branch_block_stmt_239__entry__
      -- CP-element group 0: 	 branch_block_stmt_239/$entry
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_update_start_
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_update_start_
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_update_start_
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Update/cr
      -- 
    cr_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_273_inst_req_1); -- 
    cr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_269_inst_req_1); -- 
    rr_722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => RPIPE_zeropad_input_pipe_241_inst_req_0); -- 
    cr_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_277_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_update_start_
      -- CP-element group 1: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Sample/ra
      -- 
    ra_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_241_inst_ack_0, ack => zeropad3D_CP_676_elements(1)); -- 
    cr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => RPIPE_zeropad_input_pipe_241_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_241_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Sample/$entry
      -- 
    ca_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_241_inst_ack_1, ack => zeropad3D_CP_676_elements(2)); -- 
    rr_736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => RPIPE_zeropad_input_pipe_244_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_update_start_
      -- CP-element group 3: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_sample_completed_
      -- 
    ra_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_244_inst_ack_0, ack => zeropad3D_CP_676_elements(3)); -- 
    cr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => RPIPE_zeropad_input_pipe_244_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_244_update_completed_
      -- 
    ca_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_244_inst_ack_1, ack => zeropad3D_CP_676_elements(4)); -- 
    rr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => RPIPE_zeropad_input_pipe_247_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_update_start_
      -- CP-element group 5: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Sample/ra
      -- 
    ra_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_247_inst_ack_0, ack => zeropad3D_CP_676_elements(5)); -- 
    cr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => RPIPE_zeropad_input_pipe_247_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	19 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_247_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Sample/$entry
      -- 
    ca_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_247_inst_ack_1, ack => zeropad3D_CP_676_elements(6)); -- 
    rr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_269_inst_req_0); -- 
    rr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => RPIPE_zeropad_input_pipe_250_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_update_start_
      -- CP-element group 7: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_sample_completed_
      -- 
    ra_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_250_inst_ack_0, ack => zeropad3D_CP_676_elements(7)); -- 
    cr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => RPIPE_zeropad_input_pipe_250_inst_req_1); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_250_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Sample/$entry
      -- 
    ca_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_250_inst_ack_1, ack => zeropad3D_CP_676_elements(8)); -- 
    rr_862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_273_inst_req_0); -- 
    rr_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => RPIPE_zeropad_input_pipe_253_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_update_start_
      -- CP-element group 9: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Sample/$exit
      -- 
    ra_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_253_inst_ack_0, ack => zeropad3D_CP_676_elements(9)); -- 
    cr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(9), ack => RPIPE_zeropad_input_pipe_253_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_253_Update/ca
      -- 
    ca_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_253_inst_ack_1, ack => zeropad3D_CP_676_elements(10)); -- 
    rr_876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => type_cast_277_inst_req_0); -- 
    rr_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => RPIPE_zeropad_input_pipe_256_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_update_start_
      -- 
    ra_793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_256_inst_ack_0, ack => zeropad3D_CP_676_elements(11)); -- 
    cr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(11), ack => RPIPE_zeropad_input_pipe_256_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_256_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Sample/rr
      -- 
    ca_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_256_inst_ack_1, ack => zeropad3D_CP_676_elements(12)); -- 
    rr_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(12), ack => RPIPE_zeropad_input_pipe_259_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_update_start_
      -- CP-element group 13: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Sample/$exit
      -- 
    ra_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_259_inst_ack_0, ack => zeropad3D_CP_676_elements(13)); -- 
    cr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(13), ack => RPIPE_zeropad_input_pipe_259_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_259_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Sample/rr
      -- 
    ca_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_259_inst_ack_1, ack => zeropad3D_CP_676_elements(14)); -- 
    rr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => RPIPE_zeropad_input_pipe_262_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_update_start_
      -- CP-element group 15: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Update/cr
      -- 
    ra_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_262_inst_ack_0, ack => zeropad3D_CP_676_elements(15)); -- 
    cr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(15), ack => RPIPE_zeropad_input_pipe_262_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_262_Update/$exit
      -- 
    ca_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_262_inst_ack_1, ack => zeropad3D_CP_676_elements(16)); -- 
    rr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(16), ack => RPIPE_zeropad_input_pipe_265_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_update_start_
      -- CP-element group 17: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Update/$entry
      -- 
    ra_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_265_inst_ack_0, ack => zeropad3D_CP_676_elements(17)); -- 
    cr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(17), ack => RPIPE_zeropad_input_pipe_265_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/RPIPE_zeropad_input_pipe_265_update_completed_
      -- 
    ca_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_265_inst_ack_1, ack => zeropad3D_CP_676_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	6 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Sample/$exit
      -- 
    ra_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => zeropad3D_CP_676_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_269_Update/$exit
      -- 
    ca_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => zeropad3D_CP_676_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_sample_completed_
      -- 
    ra_863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_0, ack => zeropad3D_CP_676_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_273_Update/ca
      -- 
    ca_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_1, ack => zeropad3D_CP_676_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Sample/ra
      -- 
    ra_877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_277_inst_ack_0, ack => zeropad3D_CP_676_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/type_cast_277_Update/$exit
      -- 
    ca_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_277_inst_ack_1, ack => zeropad3D_CP_676_elements(24)); -- 
    -- CP-element group 25:  branch  join  transition  place  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	22 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (10) 
      -- CP-element group 25: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300/$exit
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301__entry__
      -- CP-element group 25: 	 branch_block_stmt_239/assign_stmt_242_to_assign_stmt_300__exit__
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301_if_link/$entry
      -- CP-element group 25: 	 branch_block_stmt_239/R_cmp166_302_place
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301_eval_test/$entry
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301_eval_test/$exit
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301_eval_test/branch_req
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301_dead_link/$entry
      -- CP-element group 25: 	 branch_block_stmt_239/if_stmt_301_else_link/$entry
      -- 
    branch_req_890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(25), ack => if_stmt_301_branch_req_0); -- 
    zeropad3D_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(18) & zeropad3D_CP_676_elements(20) & zeropad3D_CP_676_elements(22) & zeropad3D_CP_676_elements(24);
      gj_zeropad3D_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  place  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	232 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_239/entry_forx_xend
      -- CP-element group 26: 	 branch_block_stmt_239/if_stmt_301_if_link/$exit
      -- CP-element group 26: 	 branch_block_stmt_239/if_stmt_301_if_link/if_choice_transition
      -- CP-element group 26: 	 branch_block_stmt_239/entry_forx_xend_PhiReq/$entry
      -- CP-element group 26: 	 branch_block_stmt_239/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_301_branch_ack_1, ack => zeropad3D_CP_676_elements(26)); -- 
    -- CP-element group 27:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	31 
    -- CP-element group 27: 	32 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (30) 
      -- CP-element group 27: 	 branch_block_stmt_239/entry_bbx_xnph
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_update_start_
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_update_start_
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348__entry__
      -- CP-element group 27: 	 branch_block_stmt_239/merge_stmt_307__exit__
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_239/if_stmt_301_else_link/else_choice_transition
      -- CP-element group 27: 	 branch_block_stmt_239/if_stmt_301_else_link/$exit
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_update_start_
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_239/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 27: 	 branch_block_stmt_239/merge_stmt_307_PhiReqMerge
      -- CP-element group 27: 	 branch_block_stmt_239/merge_stmt_307_PhiAck/$entry
      -- CP-element group 27: 	 branch_block_stmt_239/merge_stmt_307_PhiAck/$exit
      -- CP-element group 27: 	 branch_block_stmt_239/merge_stmt_307_PhiAck/dummy
      -- 
    else_choice_transition_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_301_branch_ack_0, ack => zeropad3D_CP_676_elements(27)); -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_310_inst_req_0); -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_310_inst_req_1); -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_314_inst_req_0); -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_314_inst_req_1); -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_323_inst_req_0); -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_323_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Sample/ra
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_0, ack => zeropad3D_CP_676_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_310_Update/$exit
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_1, ack => zeropad3D_CP_676_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Sample/ra
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_0, ack => zeropad3D_CP_676_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	27 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_314_Update/ca
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_1, ack => zeropad3D_CP_676_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	27 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Sample/ra
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_323_inst_ack_0, ack => zeropad3D_CP_676_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/type_cast_323_Update/ca
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_323_inst_ack_1, ack => zeropad3D_CP_676_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	226 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348/$exit
      -- CP-element group 34: 	 branch_block_stmt_239/bbx_xnph_forx_xbody
      -- CP-element group 34: 	 branch_block_stmt_239/assign_stmt_311_to_assign_stmt_348__exit__
      -- CP-element group 34: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/phi_stmt_351/$entry
      -- CP-element group 34: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/$entry
      -- 
    zeropad3D_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(29) & zeropad3D_CP_676_elements(31) & zeropad3D_CP_676_elements(33);
      gj_zeropad3D_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	231 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	74 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_sample_complete
      -- CP-element group 35: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Sample/ack
      -- 
    ack_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_offset_ack_0, ack => zeropad3D_CP_676_elements(35)); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	231 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (11) 
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_root_address_calculated
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_offset_calculated
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_base_plus_offset/$entry
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_base_plus_offset/$exit
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_base_plus_offset/sum_rename_req
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_base_plus_offset/sum_rename_ack
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_request/$entry
      -- CP-element group 36: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_request/req
      -- 
    ack_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_offset_ack_1, ack => zeropad3D_CP_676_elements(36)); -- 
    req_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(36), ack => addr_of_364_final_reg_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_request/$exit
      -- CP-element group 37: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_request/ack
      -- 
    ack_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_364_final_reg_ack_0, ack => zeropad3D_CP_676_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	231 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	71 
    -- CP-element group 38:  members (19) 
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_complete/$exit
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_complete/ack
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_word_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_root_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_address_resized
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_addr_resize/$entry
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_addr_resize/$exit
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_addr_resize/base_resize_req
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_addr_resize/base_resize_ack
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_plus_offset/$entry
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_plus_offset/$exit
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_plus_offset/sum_rename_req
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_base_plus_offset/sum_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_word_addrgen/$entry
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_word_addrgen/$exit
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_word_addrgen/root_register_req
      -- CP-element group 38: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_word_addrgen/root_register_ack
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_364_final_reg_ack_1, ack => zeropad3D_CP_676_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	231 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_update_start_
      -- CP-element group 39: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Update/cr
      -- 
    ra_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_0, ack => zeropad3D_CP_676_elements(39)); -- 
    cr_1008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(39), ack => RPIPE_zeropad_input_pipe_367_inst_req_1); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Sample/rr
      -- 
    ca_1009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_1, ack => zeropad3D_CP_676_elements(40)); -- 
    rr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => type_cast_371_inst_req_0); -- 
    rr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => RPIPE_zeropad_input_pipe_380_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Sample/ra
      -- 
    ra_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => zeropad3D_CP_676_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	231 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	71 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Update/ca
      -- 
    ca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => zeropad3D_CP_676_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	40 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_update_start_
      -- CP-element group 43: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Update/cr
      -- 
    ra_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_380_inst_ack_0, ack => zeropad3D_CP_676_elements(43)); -- 
    cr_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(43), ack => RPIPE_zeropad_input_pipe_380_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_380_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Sample/rr
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Sample/rr
      -- 
    ca_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_380_inst_ack_1, ack => zeropad3D_CP_676_elements(44)); -- 
    rr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => type_cast_384_inst_req_0); -- 
    rr_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => RPIPE_zeropad_input_pipe_398_inst_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Sample/ra
      -- 
    ra_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_384_inst_ack_0, ack => zeropad3D_CP_676_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	231 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	71 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Update/ca
      -- 
    ca_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_384_inst_ack_1, ack => zeropad3D_CP_676_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_update_start_
      -- CP-element group 47: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Update/cr
      -- 
    ra_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_398_inst_ack_0, ack => zeropad3D_CP_676_elements(47)); -- 
    cr_1064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(47), ack => RPIPE_zeropad_input_pipe_398_inst_req_1); -- 
    -- CP-element group 48:  fork  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	51 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_398_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Sample/rr
      -- 
    ca_1065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_398_inst_ack_1, ack => zeropad3D_CP_676_elements(48)); -- 
    rr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => type_cast_402_inst_req_0); -- 
    rr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => RPIPE_zeropad_input_pipe_416_inst_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Sample/ra
      -- 
    ra_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_0, ack => zeropad3D_CP_676_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	231 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	71 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Update/ca
      -- 
    ca_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_1, ack => zeropad3D_CP_676_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	48 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_update_start_
      -- CP-element group 51: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Update/cr
      -- 
    ra_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_416_inst_ack_0, ack => zeropad3D_CP_676_elements(51)); -- 
    cr_1092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(51), ack => RPIPE_zeropad_input_pipe_416_inst_req_1); -- 
    -- CP-element group 52:  fork  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (9) 
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_416_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Sample/rr
      -- 
    ca_1093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_416_inst_ack_1, ack => zeropad3D_CP_676_elements(52)); -- 
    rr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => type_cast_420_inst_req_0); -- 
    rr_1115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => RPIPE_zeropad_input_pipe_434_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Sample/ra
      -- 
    ra_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_420_inst_ack_0, ack => zeropad3D_CP_676_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	231 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	71 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Update/ca
      -- 
    ca_1107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_420_inst_ack_1, ack => zeropad3D_CP_676_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_update_start_
      -- CP-element group 55: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Update/cr
      -- 
    ra_1116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_434_inst_ack_0, ack => zeropad3D_CP_676_elements(55)); -- 
    cr_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(55), ack => RPIPE_zeropad_input_pipe_434_inst_req_1); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	59 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_434_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Sample/rr
      -- 
    ca_1121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_434_inst_ack_1, ack => zeropad3D_CP_676_elements(56)); -- 
    rr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(56), ack => type_cast_438_inst_req_0); -- 
    rr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(56), ack => RPIPE_zeropad_input_pipe_452_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Sample/ra
      -- 
    ra_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_438_inst_ack_0, ack => zeropad3D_CP_676_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	231 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	71 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Update/ca
      -- 
    ca_1135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_438_inst_ack_1, ack => zeropad3D_CP_676_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	56 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_update_start_
      -- CP-element group 59: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Update/cr
      -- 
    ra_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_452_inst_ack_0, ack => zeropad3D_CP_676_elements(59)); -- 
    cr_1148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(59), ack => RPIPE_zeropad_input_pipe_452_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	63 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_452_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Sample/rr
      -- 
    ca_1149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_452_inst_ack_1, ack => zeropad3D_CP_676_elements(60)); -- 
    rr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(60), ack => type_cast_456_inst_req_0); -- 
    rr_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(60), ack => RPIPE_zeropad_input_pipe_470_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Sample/ra
      -- 
    ra_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_0, ack => zeropad3D_CP_676_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	231 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	71 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Update/ca
      -- 
    ca_1163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_1, ack => zeropad3D_CP_676_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	60 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_update_start_
      -- CP-element group 63: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Update/cr
      -- 
    ra_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_470_inst_ack_0, ack => zeropad3D_CP_676_elements(63)); -- 
    cr_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(63), ack => RPIPE_zeropad_input_pipe_470_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	67 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_470_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Sample/rr
      -- 
    ca_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_470_inst_ack_1, ack => zeropad3D_CP_676_elements(64)); -- 
    rr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(64), ack => type_cast_474_inst_req_0); -- 
    rr_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(64), ack => RPIPE_zeropad_input_pipe_488_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Sample/ra
      -- 
    ra_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_474_inst_ack_0, ack => zeropad3D_CP_676_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	231 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	71 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Update/ca
      -- 
    ca_1191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_474_inst_ack_1, ack => zeropad3D_CP_676_elements(66)); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	64 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_update_start_
      -- CP-element group 67: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Update/cr
      -- 
    ra_1200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_488_inst_ack_0, ack => zeropad3D_CP_676_elements(67)); -- 
    cr_1204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(67), ack => RPIPE_zeropad_input_pipe_488_inst_req_1); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_488_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Sample/rr
      -- 
    ca_1205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_488_inst_ack_1, ack => zeropad3D_CP_676_elements(68)); -- 
    rr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(68), ack => type_cast_492_inst_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Sample/ra
      -- 
    ra_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_0, ack => zeropad3D_CP_676_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	231 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Update/ca
      -- 
    ca_1219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_1, ack => zeropad3D_CP_676_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	38 
    -- CP-element group 71: 	42 
    -- CP-element group 71: 	46 
    -- CP-element group 71: 	50 
    -- CP-element group 71: 	54 
    -- CP-element group 71: 	58 
    -- CP-element group 71: 	62 
    -- CP-element group 71: 	66 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/ptr_deref_500_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/ptr_deref_500_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/ptr_deref_500_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/ptr_deref_500_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/word_access_start/word_0/rr
      -- 
    rr_1257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(71), ack => ptr_deref_500_store_0_req_0); -- 
    zeropad3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(38) & zeropad3D_CP_676_elements(42) & zeropad3D_CP_676_elements(46) & zeropad3D_CP_676_elements(50) & zeropad3D_CP_676_elements(54) & zeropad3D_CP_676_elements(58) & zeropad3D_CP_676_elements(62) & zeropad3D_CP_676_elements(66) & zeropad3D_CP_676_elements(70);
      gj_zeropad3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Sample/word_access_start/word_0/ra
      -- 
    ra_1258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_500_store_0_ack_0, ack => zeropad3D_CP_676_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	231 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/word_access_complete/word_0/ca
      -- 
    ca_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_500_store_0_ack_1, ack => zeropad3D_CP_676_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	35 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514__entry__
      -- CP-element group 74: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513__exit__
      -- CP-element group 74: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/$exit
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_239/R_exitcond8_515_place
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_239/if_stmt_514_else_link/$entry
      -- 
    branch_req_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(74), ack => if_stmt_514_branch_req_0); -- 
    zeropad3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(35) & zeropad3D_CP_676_elements(73);
      gj_zeropad3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  transition  place  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	232 
    -- CP-element group 75:  members (13) 
      -- CP-element group 75: 	 branch_block_stmt_239/forx_xendx_xloopexit_forx_xend
      -- CP-element group 75: 	 branch_block_stmt_239/merge_stmt_520__exit__
      -- CP-element group 75: 	 branch_block_stmt_239/if_stmt_514_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_239/if_stmt_514_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_239/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 75: 	 branch_block_stmt_239/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_239/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_239/merge_stmt_520_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_239/merge_stmt_520_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_239/merge_stmt_520_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_239/merge_stmt_520_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_239/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_239/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_514_branch_ack_1, ack => zeropad3D_CP_676_elements(75)); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	227 
    -- CP-element group 76: 	228 
    -- CP-element group 76:  members (12) 
      -- CP-element group 76: 	 branch_block_stmt_239/if_stmt_514_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_239/if_stmt_514_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_514_branch_ack_0, ack => zeropad3D_CP_676_elements(76)); -- 
    rr_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(76), ack => type_cast_357_inst_req_0); -- 
    cr_2369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(76), ack => type_cast_357_inst_req_1); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	232 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Sample/cra
      -- 
    cra_1300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_525_call_ack_0, ack => zeropad3D_CP_676_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	232 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Update/cca
      -- CP-element group 78: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Sample/rr
      -- 
    cca_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_525_call_ack_1, ack => zeropad3D_CP_676_elements(78)); -- 
    rr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(78), ack => type_cast_530_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Sample/ra
      -- 
    ra_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_530_inst_ack_0, ack => zeropad3D_CP_676_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	232 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	193 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Update/ca
      -- 
    ca_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_530_inst_ack_1, ack => zeropad3D_CP_676_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	232 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_update_start_
      -- CP-element group 81: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Update/req
      -- 
    ack_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_532_inst_ack_0, ack => zeropad3D_CP_676_elements(81)); -- 
    req_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(81), ack => WPIPE_Block0_starting_532_inst_req_1); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Sample/req
      -- 
    ack_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_532_inst_ack_1, ack => zeropad3D_CP_676_elements(82)); -- 
    req_1341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(82), ack => WPIPE_Block0_starting_535_inst_req_0); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_update_start_
      -- CP-element group 83: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Sample/ack
      -- CP-element group 83: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Update/req
      -- 
    ack_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_535_inst_ack_0, ack => zeropad3D_CP_676_elements(83)); -- 
    req_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(83), ack => WPIPE_Block0_starting_535_inst_req_1); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_535_Update/ack
      -- CP-element group 84: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Sample/req
      -- 
    ack_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_535_inst_ack_1, ack => zeropad3D_CP_676_elements(84)); -- 
    req_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(84), ack => WPIPE_Block0_starting_538_inst_req_0); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_update_start_
      -- CP-element group 85: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Sample/ack
      -- CP-element group 85: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Update/req
      -- 
    ack_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_538_inst_ack_0, ack => zeropad3D_CP_676_elements(85)); -- 
    req_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(85), ack => WPIPE_Block0_starting_538_inst_req_1); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_538_Update/ack
      -- CP-element group 86: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Sample/req
      -- 
    ack_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_538_inst_ack_1, ack => zeropad3D_CP_676_elements(86)); -- 
    req_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(86), ack => WPIPE_Block0_starting_541_inst_req_0); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_update_start_
      -- CP-element group 87: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Update/req
      -- 
    ack_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_541_inst_ack_0, ack => zeropad3D_CP_676_elements(87)); -- 
    req_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(87), ack => WPIPE_Block0_starting_541_inst_req_1); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_541_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Sample/req
      -- 
    ack_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_541_inst_ack_1, ack => zeropad3D_CP_676_elements(88)); -- 
    req_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(88), ack => WPIPE_Block0_starting_544_inst_req_0); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_update_start_
      -- CP-element group 89: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Update/req
      -- 
    ack_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_544_inst_ack_0, ack => zeropad3D_CP_676_elements(89)); -- 
    req_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(89), ack => WPIPE_Block0_starting_544_inst_req_1); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_544_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Sample/req
      -- 
    ack_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_544_inst_ack_1, ack => zeropad3D_CP_676_elements(90)); -- 
    req_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(90), ack => WPIPE_Block0_starting_547_inst_req_0); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_update_start_
      -- CP-element group 91: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Update/req
      -- 
    ack_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_547_inst_ack_0, ack => zeropad3D_CP_676_elements(91)); -- 
    req_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(91), ack => WPIPE_Block0_starting_547_inst_req_1); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_547_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Sample/req
      -- 
    ack_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_547_inst_ack_1, ack => zeropad3D_CP_676_elements(92)); -- 
    req_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(92), ack => WPIPE_Block0_starting_550_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_update_start_
      -- CP-element group 93: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Update/req
      -- 
    ack_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_550_inst_ack_0, ack => zeropad3D_CP_676_elements(93)); -- 
    req_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(93), ack => WPIPE_Block0_starting_550_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	193 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_550_Update/ack
      -- 
    ack_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_550_inst_ack_1, ack => zeropad3D_CP_676_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	232 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_update_start_
      -- CP-element group 95: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Sample/ack
      -- CP-element group 95: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Update/req
      -- 
    ack_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_553_inst_ack_0, ack => zeropad3D_CP_676_elements(95)); -- 
    req_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(95), ack => WPIPE_Block1_starting_553_inst_req_1); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Update/ack
      -- CP-element group 96: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Sample/req
      -- 
    ack_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_553_inst_ack_1, ack => zeropad3D_CP_676_elements(96)); -- 
    req_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(96), ack => WPIPE_Block1_starting_556_inst_req_0); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Update/req
      -- CP-element group 97: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_update_start_
      -- CP-element group 97: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Sample/ack
      -- 
    ack_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_556_inst_ack_0, ack => zeropad3D_CP_676_elements(97)); -- 
    req_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(97), ack => WPIPE_Block1_starting_556_inst_req_1); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Sample/req
      -- CP-element group 98: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_Update/ack
      -- CP-element group 98: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_556_update_completed_
      -- 
    ack_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_556_inst_ack_1, ack => zeropad3D_CP_676_elements(98)); -- 
    req_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(98), ack => WPIPE_Block1_starting_559_inst_req_0); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_update_start_
      -- CP-element group 99: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Update/req
      -- 
    ack_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_559_inst_ack_0, ack => zeropad3D_CP_676_elements(99)); -- 
    req_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(99), ack => WPIPE_Block1_starting_559_inst_req_1); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Sample/req
      -- CP-element group 100: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_559_Update/$exit
      -- 
    ack_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_559_inst_ack_1, ack => zeropad3D_CP_676_elements(100)); -- 
    req_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(100), ack => WPIPE_Block1_starting_562_inst_req_0); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Update/req
      -- CP-element group 101: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_update_start_
      -- CP-element group 101: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_sample_completed_
      -- 
    ack_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_562_inst_ack_0, ack => zeropad3D_CP_676_elements(101)); -- 
    req_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(101), ack => WPIPE_Block1_starting_562_inst_req_1); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_Update/ack
      -- CP-element group 102: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_562_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Sample/req
      -- 
    ack_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_562_inst_ack_1, ack => zeropad3D_CP_676_elements(102)); -- 
    req_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(102), ack => WPIPE_Block1_starting_565_inst_req_0); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_update_start_
      -- CP-element group 103: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Update/req
      -- CP-element group 103: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Sample/ack
      -- 
    ack_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_565_inst_ack_0, ack => zeropad3D_CP_676_elements(103)); -- 
    req_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(103), ack => WPIPE_Block1_starting_565_inst_req_1); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Sample/req
      -- CP-element group 104: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_565_Update/$exit
      -- 
    ack_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_565_inst_ack_1, ack => zeropad3D_CP_676_elements(104)); -- 
    req_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(104), ack => WPIPE_Block1_starting_568_inst_req_0); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Update/req
      -- CP-element group 105: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Sample/ack
      -- CP-element group 105: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_update_start_
      -- CP-element group 105: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_sample_completed_
      -- 
    ack_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_568_inst_ack_0, ack => zeropad3D_CP_676_elements(105)); -- 
    req_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(105), ack => WPIPE_Block1_starting_568_inst_req_1); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Update/ack
      -- CP-element group 106: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Sample/req
      -- CP-element group 106: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_568_update_completed_
      -- 
    ack_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_568_inst_ack_1, ack => zeropad3D_CP_676_elements(106)); -- 
    req_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(106), ack => WPIPE_Block1_starting_571_inst_req_0); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_update_start_
      -- CP-element group 107: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Update/req
      -- CP-element group 107: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Sample/ack
      -- CP-element group 107: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Update/$entry
      -- 
    ack_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_571_inst_ack_0, ack => zeropad3D_CP_676_elements(107)); -- 
    req_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(107), ack => WPIPE_Block1_starting_571_inst_req_1); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	193 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Update/ack
      -- CP-element group 108: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_571_update_completed_
      -- 
    ack_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_571_inst_ack_1, ack => zeropad3D_CP_676_elements(108)); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	232 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_update_start_
      -- CP-element group 109: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Update/req
      -- CP-element group 109: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Sample/ack
      -- 
    ack_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_574_inst_ack_0, ack => zeropad3D_CP_676_elements(109)); -- 
    req_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(109), ack => WPIPE_Block2_starting_574_inst_req_1); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Sample/req
      -- CP-element group 110: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Update/ack
      -- CP-element group 110: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Update/$exit
      -- 
    ack_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_574_inst_ack_1, ack => zeropad3D_CP_676_elements(110)); -- 
    req_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(110), ack => WPIPE_Block2_starting_577_inst_req_0); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Update/req
      -- CP-element group 111: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Sample/ack
      -- CP-element group 111: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_update_start_
      -- 
    ack_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_577_inst_ack_0, ack => zeropad3D_CP_676_elements(111)); -- 
    req_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => WPIPE_Block2_starting_577_inst_req_1); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_577_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Sample/$entry
      -- 
    ack_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_577_inst_ack_1, ack => zeropad3D_CP_676_elements(112)); -- 
    req_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(112), ack => WPIPE_Block2_starting_580_inst_req_0); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Update/req
      -- CP-element group 113: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_update_start_
      -- 
    ack_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_580_inst_ack_0, ack => zeropad3D_CP_676_elements(113)); -- 
    req_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(113), ack => WPIPE_Block2_starting_580_inst_req_1); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Sample/req
      -- CP-element group 114: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Update/ack
      -- CP-element group 114: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_580_update_completed_
      -- 
    ack_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_580_inst_ack_1, ack => zeropad3D_CP_676_elements(114)); -- 
    req_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(114), ack => WPIPE_Block2_starting_583_inst_req_0); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Update/req
      -- CP-element group 115: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Sample/ack
      -- CP-element group 115: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_update_start_
      -- CP-element group 115: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_sample_completed_
      -- 
    ack_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_583_inst_ack_0, ack => zeropad3D_CP_676_elements(115)); -- 
    req_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(115), ack => WPIPE_Block2_starting_583_inst_req_1); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Sample/req
      -- CP-element group 116: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Update/ack
      -- CP-element group 116: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_583_update_completed_
      -- 
    ack_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_583_inst_ack_1, ack => zeropad3D_CP_676_elements(116)); -- 
    req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(116), ack => WPIPE_Block2_starting_586_inst_req_0); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (6) 
      -- CP-element group 117: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Update/req
      -- CP-element group 117: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Sample/ack
      -- CP-element group 117: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_update_start_
      -- CP-element group 117: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_sample_completed_
      -- 
    ack_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_586_inst_ack_0, ack => zeropad3D_CP_676_elements(117)); -- 
    req_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(117), ack => WPIPE_Block2_starting_586_inst_req_1); -- 
    -- CP-element group 118:  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (6) 
      -- CP-element group 118: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Sample/req
      -- CP-element group 118: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Update/ack
      -- CP-element group 118: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_586_update_completed_
      -- 
    ack_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_586_inst_ack_1, ack => zeropad3D_CP_676_elements(118)); -- 
    req_1593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(118), ack => WPIPE_Block2_starting_589_inst_req_0); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Update/req
      -- CP-element group 119: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Sample/ack
      -- CP-element group 119: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_update_start_
      -- CP-element group 119: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_sample_completed_
      -- 
    ack_1594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_589_inst_ack_0, ack => zeropad3D_CP_676_elements(119)); -- 
    req_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(119), ack => WPIPE_Block2_starting_589_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Update/ack
      -- CP-element group 120: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Sample/req
      -- CP-element group 120: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_589_update_completed_
      -- 
    ack_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_589_inst_ack_1, ack => zeropad3D_CP_676_elements(120)); -- 
    req_1607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(120), ack => WPIPE_Block2_starting_592_inst_req_0); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Update/req
      -- CP-element group 121: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_update_start_
      -- CP-element group 121: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Sample/$exit
      -- 
    ack_1608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_592_inst_ack_0, ack => zeropad3D_CP_676_elements(121)); -- 
    req_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(121), ack => WPIPE_Block2_starting_592_inst_req_1); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	193 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_Update/ack
      -- CP-element group 122: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_592_update_completed_
      -- 
    ack_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_592_inst_ack_1, ack => zeropad3D_CP_676_elements(122)); -- 
    -- CP-element group 123:  transition  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	232 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (6) 
      -- CP-element group 123: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Sample/ack
      -- CP-element group 123: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Update/req
      -- CP-element group 123: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_update_start_
      -- 
    ack_1622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_595_inst_ack_0, ack => zeropad3D_CP_676_elements(123)); -- 
    req_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(123), ack => WPIPE_Block3_starting_595_inst_req_1); -- 
    -- CP-element group 124:  transition  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Update/ack
      -- CP-element group 124: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Sample/req
      -- CP-element group 124: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Sample/$entry
      -- 
    ack_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_595_inst_ack_1, ack => zeropad3D_CP_676_elements(124)); -- 
    req_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => WPIPE_Block3_starting_598_inst_req_0); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (6) 
      -- CP-element group 125: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Update/req
      -- CP-element group 125: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_update_start_
      -- 
    ack_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_598_inst_ack_0, ack => zeropad3D_CP_676_elements(125)); -- 
    req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(125), ack => WPIPE_Block3_starting_598_inst_req_1); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Sample/req
      -- CP-element group 126: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_598_update_completed_
      -- 
    ack_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_598_inst_ack_1, ack => zeropad3D_CP_676_elements(126)); -- 
    req_1649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(126), ack => WPIPE_Block3_starting_601_inst_req_0); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (6) 
      -- CP-element group 127: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Update/req
      -- CP-element group 127: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Sample/ack
      -- CP-element group 127: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_update_start_
      -- CP-element group 127: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Update/$entry
      -- 
    ack_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_601_inst_ack_0, ack => zeropad3D_CP_676_elements(127)); -- 
    req_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(127), ack => WPIPE_Block3_starting_601_inst_req_1); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_Update/ack
      -- CP-element group 128: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Sample/req
      -- CP-element group 128: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_601_update_completed_
      -- 
    ack_1655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_601_inst_ack_1, ack => zeropad3D_CP_676_elements(128)); -- 
    req_1663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => WPIPE_Block3_starting_604_inst_req_0); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_update_start_
      -- CP-element group 129: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Sample/ack
      -- CP-element group 129: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Update/req
      -- 
    ack_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_604_inst_ack_0, ack => zeropad3D_CP_676_elements(129)); -- 
    req_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(129), ack => WPIPE_Block3_starting_604_inst_req_1); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Sample/req
      -- CP-element group 130: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_604_Update/ack
      -- 
    ack_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_604_inst_ack_1, ack => zeropad3D_CP_676_elements(130)); -- 
    req_1677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(130), ack => WPIPE_Block3_starting_607_inst_req_0); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Update/req
      -- CP-element group 131: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Sample/ack
      -- CP-element group 131: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_update_start_
      -- CP-element group 131: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_sample_completed_
      -- 
    ack_1678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_607_inst_ack_0, ack => zeropad3D_CP_676_elements(131)); -- 
    req_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(131), ack => WPIPE_Block3_starting_607_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Sample/req
      -- CP-element group 132: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_607_update_completed_
      -- 
    ack_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_607_inst_ack_1, ack => zeropad3D_CP_676_elements(132)); -- 
    req_1691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(132), ack => WPIPE_Block3_starting_610_inst_req_0); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Update/req
      -- CP-element group 133: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Sample/ack
      -- CP-element group 133: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_update_start_
      -- CP-element group 133: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_sample_completed_
      -- 
    ack_1692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_610_inst_ack_0, ack => zeropad3D_CP_676_elements(133)); -- 
    req_1696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(133), ack => WPIPE_Block3_starting_610_inst_req_1); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Sample/req
      -- CP-element group 134: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Update/ack
      -- CP-element group 134: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_610_update_completed_
      -- 
    ack_1697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_610_inst_ack_1, ack => zeropad3D_CP_676_elements(134)); -- 
    req_1705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(134), ack => WPIPE_Block3_starting_613_inst_req_0); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_update_start_
      -- CP-element group 135: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Update/req
      -- CP-element group 135: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Sample/ack
      -- 
    ack_1706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_613_inst_ack_0, ack => zeropad3D_CP_676_elements(135)); -- 
    req_1710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(135), ack => WPIPE_Block3_starting_613_inst_req_1); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	193 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Update/ack
      -- CP-element group 136: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_613_Update/$exit
      -- 
    ack_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_613_inst_ack_1, ack => zeropad3D_CP_676_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	232 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Update/req
      -- CP-element group 137: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_update_start_
      -- CP-element group 137: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_sample_completed_
      -- 
    ack_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_616_inst_ack_0, ack => zeropad3D_CP_676_elements(137)); -- 
    req_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(137), ack => WPIPE_Block4_starting_616_inst_req_1); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Sample/req
      -- CP-element group 138: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Update/ack
      -- CP-element group 138: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_update_completed_
      -- 
    ack_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_616_inst_ack_1, ack => zeropad3D_CP_676_elements(138)); -- 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(138), ack => WPIPE_Block4_starting_619_inst_req_0); -- 
    -- CP-element group 139:  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (6) 
      -- CP-element group 139: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_update_start_
      -- CP-element group 139: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Sample/ack
      -- CP-element group 139: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Update/req
      -- 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_619_inst_ack_0, ack => zeropad3D_CP_676_elements(139)); -- 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(139), ack => WPIPE_Block4_starting_619_inst_req_1); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Sample/req
      -- CP-element group 140: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_619_Update/ack
      -- 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_619_inst_ack_1, ack => zeropad3D_CP_676_elements(140)); -- 
    req_1747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(140), ack => WPIPE_Block4_starting_622_inst_req_0); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Update/req
      -- CP-element group 141: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Sample/ack
      -- CP-element group 141: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_update_start_
      -- CP-element group 141: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_sample_completed_
      -- 
    ack_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_622_inst_ack_0, ack => zeropad3D_CP_676_elements(141)); -- 
    req_1752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(141), ack => WPIPE_Block4_starting_622_inst_req_1); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Update/ack
      -- CP-element group 142: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Sample/req
      -- CP-element group 142: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_622_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_sample_start_
      -- 
    ack_1753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_622_inst_ack_1, ack => zeropad3D_CP_676_elements(142)); -- 
    req_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(142), ack => WPIPE_Block4_starting_625_inst_req_0); -- 
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (6) 
      -- CP-element group 143: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Sample/ack
      -- CP-element group 143: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_update_start_
      -- CP-element group 143: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Update/req
      -- CP-element group 143: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Update/$entry
      -- 
    ack_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_625_inst_ack_0, ack => zeropad3D_CP_676_elements(143)); -- 
    req_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(143), ack => WPIPE_Block4_starting_625_inst_req_1); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Sample/req
      -- CP-element group 144: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Update/ack
      -- CP-element group 144: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_625_Update/$exit
      -- 
    ack_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_625_inst_ack_1, ack => zeropad3D_CP_676_elements(144)); -- 
    req_1775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(144), ack => WPIPE_Block4_starting_628_inst_req_0); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Sample/ack
      -- CP-element group 145: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Update/req
      -- CP-element group 145: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_update_start_
      -- CP-element group 145: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_sample_completed_
      -- 
    ack_1776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_628_inst_ack_0, ack => zeropad3D_CP_676_elements(145)); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(145), ack => WPIPE_Block4_starting_628_inst_req_1); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Update/ack
      -- CP-element group 146: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_628_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Sample/req
      -- CP-element group 146: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Sample/$entry
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_628_inst_ack_1, ack => zeropad3D_CP_676_elements(146)); -- 
    req_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(146), ack => WPIPE_Block4_starting_631_inst_req_0); -- 
    -- CP-element group 147:  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Update/req
      -- CP-element group 147: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Sample/ack
      -- CP-element group 147: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_update_start_
      -- 
    ack_1790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_631_inst_ack_0, ack => zeropad3D_CP_676_elements(147)); -- 
    req_1794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(147), ack => WPIPE_Block4_starting_631_inst_req_1); -- 
    -- CP-element group 148:  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Sample/req
      -- CP-element group 148: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Update/ack
      -- CP-element group 148: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_631_update_completed_
      -- 
    ack_1795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_631_inst_ack_1, ack => zeropad3D_CP_676_elements(148)); -- 
    req_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(148), ack => WPIPE_Block4_starting_634_inst_req_0); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Sample/ack
      -- CP-element group 149: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Update/req
      -- CP-element group 149: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_update_start_
      -- CP-element group 149: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_sample_completed_
      -- 
    ack_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_634_inst_ack_0, ack => zeropad3D_CP_676_elements(149)); -- 
    req_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => WPIPE_Block4_starting_634_inst_req_1); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	193 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_Update/ack
      -- CP-element group 150: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_634_update_completed_
      -- 
    ack_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_starting_634_inst_ack_1, ack => zeropad3D_CP_676_elements(150)); -- 
    -- CP-element group 151:  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	232 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (6) 
      -- CP-element group 151: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Update/req
      -- CP-element group 151: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Sample/ack
      -- CP-element group 151: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_update_start_
      -- 
    ack_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_637_inst_ack_0, ack => zeropad3D_CP_676_elements(151)); -- 
    req_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => WPIPE_Block5_starting_637_inst_req_1); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Sample/req
      -- CP-element group 152: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_update_completed_
      -- 
    ack_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_637_inst_ack_1, ack => zeropad3D_CP_676_elements(152)); -- 
    req_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(152), ack => WPIPE_Block5_starting_640_inst_req_0); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Sample/ack
      -- CP-element group 153: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Update/req
      -- CP-element group 153: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_update_start_
      -- 
    ack_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_640_inst_ack_0, ack => zeropad3D_CP_676_elements(153)); -- 
    req_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(153), ack => WPIPE_Block5_starting_640_inst_req_1); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Update/ack
      -- CP-element group 154: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_640_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Sample/req
      -- 
    ack_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_640_inst_ack_1, ack => zeropad3D_CP_676_elements(154)); -- 
    req_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(154), ack => WPIPE_Block5_starting_643_inst_req_0); -- 
    -- CP-element group 155:  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_update_start_
      -- CP-element group 155: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Update/req
      -- CP-element group 155: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Sample/ack
      -- 
    ack_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_643_inst_ack_0, ack => zeropad3D_CP_676_elements(155)); -- 
    req_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(155), ack => WPIPE_Block5_starting_643_inst_req_1); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Sample/req
      -- CP-element group 156: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_643_Update/$exit
      -- 
    ack_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_643_inst_ack_1, ack => zeropad3D_CP_676_elements(156)); -- 
    req_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(156), ack => WPIPE_Block5_starting_646_inst_req_0); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Update/req
      -- CP-element group 157: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Sample/ack
      -- CP-element group 157: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_update_start_
      -- CP-element group 157: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_sample_completed_
      -- 
    ack_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_646_inst_ack_0, ack => zeropad3D_CP_676_elements(157)); -- 
    req_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => WPIPE_Block5_starting_646_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Update/ack
      -- CP-element group 158: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Sample/req
      -- CP-element group 158: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_646_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_sample_start_
      -- 
    ack_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_646_inst_ack_1, ack => zeropad3D_CP_676_elements(158)); -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(158), ack => WPIPE_Block5_starting_649_inst_req_0); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Sample/ack
      -- CP-element group 159: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_update_start_
      -- CP-element group 159: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Update/req
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_649_inst_ack_0, ack => zeropad3D_CP_676_elements(159)); -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(159), ack => WPIPE_Block5_starting_649_inst_req_1); -- 
    -- CP-element group 160:  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Update/ack
      -- CP-element group 160: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Sample/req
      -- CP-element group 160: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_649_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Sample/$entry
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_649_inst_ack_1, ack => zeropad3D_CP_676_elements(160)); -- 
    req_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(160), ack => WPIPE_Block5_starting_652_inst_req_0); -- 
    -- CP-element group 161:  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (6) 
      -- CP-element group 161: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_update_start_
      -- CP-element group 161: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Update/req
      -- CP-element group 161: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Sample/ack
      -- 
    ack_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_652_inst_ack_0, ack => zeropad3D_CP_676_elements(161)); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(161), ack => WPIPE_Block5_starting_652_inst_req_1); -- 
    -- CP-element group 162:  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (6) 
      -- CP-element group 162: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Update/ack
      -- CP-element group 162: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Sample/req
      -- CP-element group 162: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_652_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Sample/$entry
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_652_inst_ack_1, ack => zeropad3D_CP_676_elements(162)); -- 
    req_1901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(162), ack => WPIPE_Block5_starting_655_inst_req_0); -- 
    -- CP-element group 163:  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Update/req
      -- CP-element group 163: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Sample/ack
      -- CP-element group 163: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_update_start_
      -- 
    ack_1902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_655_inst_ack_0, ack => zeropad3D_CP_676_elements(163)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(163), ack => WPIPE_Block5_starting_655_inst_req_1); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	193 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Update/ack
      -- CP-element group 164: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_655_update_completed_
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_starting_655_inst_ack_1, ack => zeropad3D_CP_676_elements(164)); -- 
    -- CP-element group 165:  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	232 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (6) 
      -- CP-element group 165: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_update_start_
      -- CP-element group 165: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Sample/ack
      -- CP-element group 165: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Update/req
      -- 
    ack_1916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_658_inst_ack_0, ack => zeropad3D_CP_676_elements(165)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(165), ack => WPIPE_Block6_starting_658_inst_req_1); -- 
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Update/ack
      -- CP-element group 166: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Sample/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_658_inst_ack_1, ack => zeropad3D_CP_676_elements(166)); -- 
    req_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => WPIPE_Block6_starting_661_inst_req_0); -- 
    -- CP-element group 167:  transition  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167:  members (6) 
      -- CP-element group 167: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_update_start_
      -- CP-element group 167: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Sample/ack
      -- CP-element group 167: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Update/req
      -- 
    ack_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_661_inst_ack_0, ack => zeropad3D_CP_676_elements(167)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => WPIPE_Block6_starting_661_inst_req_1); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_661_Update/ack
      -- CP-element group 168: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Sample/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_661_inst_ack_1, ack => zeropad3D_CP_676_elements(168)); -- 
    req_1943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(168), ack => WPIPE_Block6_starting_664_inst_req_0); -- 
    -- CP-element group 169:  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (6) 
      -- CP-element group 169: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_update_start_
      -- CP-element group 169: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Update/req
      -- 
    ack_1944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_664_inst_ack_0, ack => zeropad3D_CP_676_elements(169)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(169), ack => WPIPE_Block6_starting_664_inst_req_1); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_664_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Sample/req
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_664_inst_ack_1, ack => zeropad3D_CP_676_elements(170)); -- 
    req_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(170), ack => WPIPE_Block6_starting_667_inst_req_0); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_update_start_
      -- CP-element group 171: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Update/req
      -- 
    ack_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_667_inst_ack_0, ack => zeropad3D_CP_676_elements(171)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(171), ack => WPIPE_Block6_starting_667_inst_req_1); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_667_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Sample/req
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_667_inst_ack_1, ack => zeropad3D_CP_676_elements(172)); -- 
    req_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => WPIPE_Block6_starting_670_inst_req_0); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_update_start_
      -- CP-element group 173: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Sample/ack
      -- CP-element group 173: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Update/req
      -- 
    ack_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_670_inst_ack_0, ack => zeropad3D_CP_676_elements(173)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(173), ack => WPIPE_Block6_starting_670_inst_req_1); -- 
    -- CP-element group 174:  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (6) 
      -- CP-element group 174: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_670_Update/ack
      -- CP-element group 174: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Sample/req
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_670_inst_ack_1, ack => zeropad3D_CP_676_elements(174)); -- 
    req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(174), ack => WPIPE_Block6_starting_673_inst_req_0); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_update_start_
      -- CP-element group 175: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Sample/ack
      -- CP-element group 175: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Update/req
      -- 
    ack_1986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_673_inst_ack_0, ack => zeropad3D_CP_676_elements(175)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => WPIPE_Block6_starting_673_inst_req_1); -- 
    -- CP-element group 176:  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (6) 
      -- CP-element group 176: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_673_Update/ack
      -- CP-element group 176: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Sample/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_673_inst_ack_1, ack => zeropad3D_CP_676_elements(176)); -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(176), ack => WPIPE_Block6_starting_676_inst_req_0); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_update_start_
      -- CP-element group 177: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Sample/ack
      -- CP-element group 177: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Update/req
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_676_inst_ack_0, ack => zeropad3D_CP_676_elements(177)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(177), ack => WPIPE_Block6_starting_676_inst_req_1); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	193 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_676_Update/ack
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_starting_676_inst_ack_1, ack => zeropad3D_CP_676_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	232 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_update_start_
      -- CP-element group 179: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Sample/ack
      -- CP-element group 179: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Update/req
      -- 
    ack_2014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_679_inst_ack_0, ack => zeropad3D_CP_676_elements(179)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(179), ack => WPIPE_Block7_starting_679_inst_req_1); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Update/ack
      -- CP-element group 180: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Sample/req
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_679_inst_ack_1, ack => zeropad3D_CP_676_elements(180)); -- 
    req_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(180), ack => WPIPE_Block7_starting_682_inst_req_0); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_update_start_
      -- CP-element group 181: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Sample/ack
      -- CP-element group 181: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Update/req
      -- 
    ack_2028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_682_inst_ack_0, ack => zeropad3D_CP_676_elements(181)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(181), ack => WPIPE_Block7_starting_682_inst_req_1); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_682_Update/ack
      -- CP-element group 182: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Sample/req
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_682_inst_ack_1, ack => zeropad3D_CP_676_elements(182)); -- 
    req_2041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(182), ack => WPIPE_Block7_starting_685_inst_req_0); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_update_start_
      -- CP-element group 183: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Sample/ack
      -- CP-element group 183: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Update/req
      -- 
    ack_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_685_inst_ack_0, ack => zeropad3D_CP_676_elements(183)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(183), ack => WPIPE_Block7_starting_685_inst_req_1); -- 
    -- CP-element group 184:  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (6) 
      -- CP-element group 184: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_685_Update/ack
      -- CP-element group 184: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Sample/req
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_685_inst_ack_1, ack => zeropad3D_CP_676_elements(184)); -- 
    req_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(184), ack => WPIPE_Block7_starting_688_inst_req_0); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_update_start_
      -- CP-element group 185: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Sample/ack
      -- CP-element group 185: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Update/req
      -- 
    ack_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_688_inst_ack_0, ack => zeropad3D_CP_676_elements(185)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(185), ack => WPIPE_Block7_starting_688_inst_req_1); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_688_Update/ack
      -- CP-element group 186: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Sample/req
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_688_inst_ack_1, ack => zeropad3D_CP_676_elements(186)); -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(186), ack => WPIPE_Block7_starting_691_inst_req_0); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_update_start_
      -- CP-element group 187: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Update/req
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_691_inst_ack_0, ack => zeropad3D_CP_676_elements(187)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(187), ack => WPIPE_Block7_starting_691_inst_req_1); -- 
    -- CP-element group 188:  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (6) 
      -- CP-element group 188: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_691_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Sample/req
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_691_inst_ack_1, ack => zeropad3D_CP_676_elements(188)); -- 
    req_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(188), ack => WPIPE_Block7_starting_694_inst_req_0); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_update_start_
      -- CP-element group 189: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Sample/ack
      -- CP-element group 189: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Update/req
      -- 
    ack_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_694_inst_ack_0, ack => zeropad3D_CP_676_elements(189)); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(189), ack => WPIPE_Block7_starting_694_inst_req_1); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_694_Update/ack
      -- CP-element group 190: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Sample/req
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_694_inst_ack_1, ack => zeropad3D_CP_676_elements(190)); -- 
    req_2097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(190), ack => WPIPE_Block7_starting_697_inst_req_0); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_update_start_
      -- CP-element group 191: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Sample/ack
      -- CP-element group 191: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Update/req
      -- 
    ack_2098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_697_inst_ack_0, ack => zeropad3D_CP_676_elements(191)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(191), ack => WPIPE_Block7_starting_697_inst_req_1); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_697_Update/ack
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_starting_697_inst_ack_1, ack => zeropad3D_CP_676_elements(192)); -- 
    -- CP-element group 193:  join  fork  transition  place  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	80 
    -- CP-element group 193: 	94 
    -- CP-element group 193: 	108 
    -- CP-element group 193: 	122 
    -- CP-element group 193: 	136 
    -- CP-element group 193: 	150 
    -- CP-element group 193: 	164 
    -- CP-element group 193: 	178 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193: 	196 
    -- CP-element group 193: 	198 
    -- CP-element group 193: 	200 
    -- CP-element group 193: 	202 
    -- CP-element group 193: 	204 
    -- CP-element group 193: 	206 
    -- CP-element group 193: 	208 
    -- CP-element group 193:  members (28) 
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724__entry__
      -- CP-element group 193: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699__exit__
      -- CP-element group 193: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/$exit
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Sample/rr
      -- 
    rr_2114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block0_complete_702_inst_req_0); -- 
    rr_2128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block1_complete_705_inst_req_0); -- 
    rr_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block2_complete_708_inst_req_0); -- 
    rr_2156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block3_complete_711_inst_req_0); -- 
    rr_2170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block4_complete_714_inst_req_0); -- 
    rr_2184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block5_complete_717_inst_req_0); -- 
    rr_2198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block6_complete_720_inst_req_0); -- 
    rr_2212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => RPIPE_Block7_complete_723_inst_req_0); -- 
    zeropad3D_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(80) & zeropad3D_CP_676_elements(94) & zeropad3D_CP_676_elements(108) & zeropad3D_CP_676_elements(122) & zeropad3D_CP_676_elements(136) & zeropad3D_CP_676_elements(150) & zeropad3D_CP_676_elements(164) & zeropad3D_CP_676_elements(178) & zeropad3D_CP_676_elements(192);
      gj_zeropad3D_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_update_start_
      -- CP-element group 194: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Update/cr
      -- 
    ra_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_702_inst_ack_0, ack => zeropad3D_CP_676_elements(194)); -- 
    cr_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(194), ack => RPIPE_Block0_complete_702_inst_req_1); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	210 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block0_complete_702_Update/ca
      -- 
    ca_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_702_inst_ack_1, ack => zeropad3D_CP_676_elements(195)); -- 
    -- CP-element group 196:  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	193 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (6) 
      -- CP-element group 196: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_update_start_
      -- CP-element group 196: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Sample/ra
      -- CP-element group 196: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Update/$entry
      -- CP-element group 196: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Update/cr
      -- 
    ra_2129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_complete_705_inst_ack_0, ack => zeropad3D_CP_676_elements(196)); -- 
    cr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(196), ack => RPIPE_Block1_complete_705_inst_req_1); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	210 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block1_complete_705_Update/ca
      -- 
    ca_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_complete_705_inst_ack_1, ack => zeropad3D_CP_676_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	193 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_update_start_
      -- CP-element group 198: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Update/cr
      -- 
    ra_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_complete_708_inst_ack_0, ack => zeropad3D_CP_676_elements(198)); -- 
    cr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(198), ack => RPIPE_Block2_complete_708_inst_req_1); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	210 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block2_complete_708_Update/ca
      -- 
    ca_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_complete_708_inst_ack_1, ack => zeropad3D_CP_676_elements(199)); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	193 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_update_start_
      -- CP-element group 200: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Update/cr
      -- 
    ra_2157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_complete_711_inst_ack_0, ack => zeropad3D_CP_676_elements(200)); -- 
    cr_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(200), ack => RPIPE_Block3_complete_711_inst_req_1); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	210 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block3_complete_711_Update/ca
      -- 
    ca_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_complete_711_inst_ack_1, ack => zeropad3D_CP_676_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	193 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_update_start_
      -- CP-element group 202: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Update/cr
      -- 
    ra_2171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_complete_714_inst_ack_0, ack => zeropad3D_CP_676_elements(202)); -- 
    cr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(202), ack => RPIPE_Block4_complete_714_inst_req_1); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	210 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block4_complete_714_Update/ca
      -- 
    ca_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_complete_714_inst_ack_1, ack => zeropad3D_CP_676_elements(203)); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	193 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_update_start_
      -- CP-element group 204: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Update/cr
      -- 
    ra_2185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_complete_717_inst_ack_0, ack => zeropad3D_CP_676_elements(204)); -- 
    cr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(204), ack => RPIPE_Block5_complete_717_inst_req_1); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	210 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block5_complete_717_Update/ca
      -- 
    ca_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_complete_717_inst_ack_1, ack => zeropad3D_CP_676_elements(205)); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	193 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_update_start_
      -- CP-element group 206: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Sample/ra
      -- CP-element group 206: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Update/cr
      -- 
    ra_2199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_complete_720_inst_ack_0, ack => zeropad3D_CP_676_elements(206)); -- 
    cr_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(206), ack => RPIPE_Block6_complete_720_inst_req_1); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	210 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block6_complete_720_Update/ca
      -- 
    ca_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_complete_720_inst_ack_1, ack => zeropad3D_CP_676_elements(207)); -- 
    -- CP-element group 208:  transition  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	193 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_update_start_
      -- CP-element group 208: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Sample/ra
      -- CP-element group 208: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Update/cr
      -- 
    ra_2213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_complete_723_inst_ack_0, ack => zeropad3D_CP_676_elements(208)); -- 
    cr_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(208), ack => RPIPE_Block7_complete_723_inst_req_1); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/RPIPE_Block7_complete_723_Update/ca
      -- 
    ca_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_complete_723_inst_ack_1, ack => zeropad3D_CP_676_elements(209)); -- 
    -- CP-element group 210:  join  fork  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	195 
    -- CP-element group 210: 	197 
    -- CP-element group 210: 	199 
    -- CP-element group 210: 	201 
    -- CP-element group 210: 	203 
    -- CP-element group 210: 	205 
    -- CP-element group 210: 	207 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210: 	214 
    -- CP-element group 210:  members (13) 
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740__entry__
      -- CP-element group 210: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724__exit__
      -- CP-element group 210: 	 branch_block_stmt_239/assign_stmt_703_to_assign_stmt_724/$exit
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/$entry
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_update_start_
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Sample/crr
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Update/ccr
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_update_start_
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Update/cr
      -- 
    crr_2229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => call_stmt_727_call_req_0); -- 
    ccr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => call_stmt_727_call_req_1); -- 
    cr_2248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_731_inst_req_1); -- 
    zeropad3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(195) & zeropad3D_CP_676_elements(197) & zeropad3D_CP_676_elements(199) & zeropad3D_CP_676_elements(201) & zeropad3D_CP_676_elements(203) & zeropad3D_CP_676_elements(205) & zeropad3D_CP_676_elements(207) & zeropad3D_CP_676_elements(209);
      gj_zeropad3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Sample/cra
      -- 
    cra_2230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_727_call_ack_0, ack => zeropad3D_CP_676_elements(211)); -- 
    -- CP-element group 212:  transition  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (6) 
      -- CP-element group 212: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/call_stmt_727_Update/cca
      -- CP-element group 212: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Sample/rr
      -- 
    cca_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_727_call_ack_1, ack => zeropad3D_CP_676_elements(212)); -- 
    rr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(212), ack => type_cast_731_inst_req_0); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Sample/ra
      -- 
    ra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => zeropad3D_CP_676_elements(213)); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	210 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/type_cast_731_Update/ca
      -- CP-element group 214: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Sample/req
      -- 
    ca_2249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => zeropad3D_CP_676_elements(214)); -- 
    req_2257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(214), ack => WPIPE_elapsed_time_pipe_738_inst_req_0); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_update_start_
      -- CP-element group 215: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Update/req
      -- 
    ack_2258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_738_inst_ack_0, ack => zeropad3D_CP_676_elements(215)); -- 
    req_2262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(215), ack => WPIPE_elapsed_time_pipe_738_inst_req_1); -- 
    -- CP-element group 216:  fork  transition  place  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216: 	218 
    -- CP-element group 216: 	219 
    -- CP-element group 216: 	220 
    -- CP-element group 216: 	221 
    -- CP-element group 216: 	222 
    -- CP-element group 216: 	225 
    -- CP-element group 216:  members (28) 
      -- CP-element group 216: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740__exit__
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765__entry__
      -- CP-element group 216: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/$exit
      -- CP-element group 216: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_239/call_stmt_727_to_assign_stmt_740/WPIPE_elapsed_time_pipe_738_Update/ack
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_update_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Sample/rr
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Update/cr
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_update_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Sample/rr
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Update/cr
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_update_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Sample/rr
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Update/cr
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_update_start_
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Update/ccr
      -- 
    ack_2263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_738_inst_ack_1, ack => zeropad3D_CP_676_elements(216)); -- 
    rr_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => type_cast_744_inst_req_0); -- 
    cr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => type_cast_744_inst_req_1); -- 
    rr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => type_cast_748_inst_req_0); -- 
    cr_2293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => type_cast_748_inst_req_1); -- 
    rr_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => type_cast_752_inst_req_0); -- 
    cr_2307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => type_cast_752_inst_req_1); -- 
    ccr_2321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(216), ack => call_stmt_765_call_req_1); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Sample/ra
      -- 
    ra_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_744_inst_ack_0, ack => zeropad3D_CP_676_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	223 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_744_Update/ca
      -- 
    ca_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_744_inst_ack_1, ack => zeropad3D_CP_676_elements(218)); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	216 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Sample/ra
      -- 
    ra_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_748_inst_ack_0, ack => zeropad3D_CP_676_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	216 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_748_Update/ca
      -- 
    ca_2294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_748_inst_ack_1, ack => zeropad3D_CP_676_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	216 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Sample/ra
      -- 
    ra_2303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_0, ack => zeropad3D_CP_676_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	216 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/type_cast_752_Update/ca
      -- 
    ca_2308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_1, ack => zeropad3D_CP_676_elements(222)); -- 
    -- CP-element group 223:  join  transition  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	218 
    -- CP-element group 223: 	220 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Sample/crr
      -- 
    crr_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(223), ack => call_stmt_765_call_req_0); -- 
    zeropad3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(218) & zeropad3D_CP_676_elements(220) & zeropad3D_CP_676_elements(222);
      gj_zeropad3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Sample/cra
      -- 
    cra_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_765_call_ack_0, ack => zeropad3D_CP_676_elements(224)); -- 
    -- CP-element group 225:  transition  place  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	216 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (16) 
      -- CP-element group 225: 	 $exit
      -- CP-element group 225: 	 branch_block_stmt_239/merge_stmt_767_PhiAck/$exit
      -- CP-element group 225: 	 branch_block_stmt_239/return__
      -- CP-element group 225: 	 branch_block_stmt_239/branch_block_stmt_239__exit__
      -- CP-element group 225: 	 branch_block_stmt_239/merge_stmt_767__exit__
      -- CP-element group 225: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765__exit__
      -- CP-element group 225: 	 branch_block_stmt_239/$exit
      -- CP-element group 225: 	 branch_block_stmt_239/merge_stmt_767_PhiAck/dummy
      -- CP-element group 225: 	 branch_block_stmt_239/return___PhiReq/$exit
      -- CP-element group 225: 	 branch_block_stmt_239/merge_stmt_767_PhiAck/$entry
      -- CP-element group 225: 	 branch_block_stmt_239/return___PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/$exit
      -- CP-element group 225: 	 branch_block_stmt_239/merge_stmt_767_PhiReqMerge
      -- CP-element group 225: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_239/assign_stmt_745_to_call_stmt_765/call_stmt_765_Update/cca
      -- 
    cca_2322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_765_call_ack_1, ack => zeropad3D_CP_676_elements(225)); -- 
    -- CP-element group 226:  transition  output  delay-element  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	34 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	230 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 226: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/phi_stmt_351/$exit
      -- CP-element group 226: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/$exit
      -- CP-element group 226: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_355_konst_delay_trans
      -- CP-element group 226: 	 branch_block_stmt_239/bbx_xnph_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_req
      -- 
    phi_stmt_351_req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_351_req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(226), ack => phi_stmt_351_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(226) is a control-delay.
    cp_element_226_delay: control_delay_element  generic map(name => " 226_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(34), ack => zeropad3D_CP_676_elements(226), clk => clk, reset =>reset);
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	76 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (2) 
      -- CP-element group 227: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Sample/ra
      -- 
    ra_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => zeropad3D_CP_676_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	76 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/Update/ca
      -- 
    ca_2370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => zeropad3D_CP_676_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (6) 
      -- CP-element group 229: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/$exit
      -- CP-element group 229: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/$exit
      -- CP-element group 229: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/$exit
      -- CP-element group 229: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_sources/type_cast_357/SplitProtocol/$exit
      -- CP-element group 229: 	 branch_block_stmt_239/forx_xbody_forx_xbody_PhiReq/phi_stmt_351/phi_stmt_351_req
      -- 
    phi_stmt_351_req_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_351_req_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(229), ack => phi_stmt_351_req_1); -- 
    zeropad3D_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(227) & zeropad3D_CP_676_elements(228);
      gj_zeropad3D_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  merge  transition  place  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	226 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (2) 
      -- CP-element group 230: 	 branch_block_stmt_239/merge_stmt_350_PhiReqMerge
      -- CP-element group 230: 	 branch_block_stmt_239/merge_stmt_350_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(230) <= OrReduce(zeropad3D_CP_676_elements(226) & zeropad3D_CP_676_elements(229));
    -- CP-element group 231:  fork  transition  place  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	35 
    -- CP-element group 231: 	36 
    -- CP-element group 231: 	38 
    -- CP-element group 231: 	39 
    -- CP-element group 231: 	42 
    -- CP-element group 231: 	46 
    -- CP-element group 231: 	50 
    -- CP-element group 231: 	54 
    -- CP-element group 231: 	58 
    -- CP-element group 231: 	62 
    -- CP-element group 231: 	66 
    -- CP-element group 231: 	70 
    -- CP-element group 231: 	73 
    -- CP-element group 231:  members (56) 
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513__entry__
      -- CP-element group 231: 	 branch_block_stmt_239/merge_stmt_350__exit__
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_resized_1
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_scaled_1
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_computed_1
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_resize_1/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_resize_1/$exit
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_resize_1/index_resize_req
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_resize_1/index_resize_ack
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_scale_1/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_scale_1/$exit
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_scale_1/scale_rename_req
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_index_scale_1/scale_rename_ack
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_update_start
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Sample/req
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/array_obj_ref_363_final_index_sum_regn_Update/req
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_complete/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/addr_of_364_complete/req
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/RPIPE_zeropad_input_pipe_367_Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_371_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_384_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_402_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_420_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_438_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_456_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_474_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/type_cast_492_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_update_start_
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/word_access_complete/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/word_access_complete/word_0/$entry
      -- CP-element group 231: 	 branch_block_stmt_239/assign_stmt_365_to_assign_stmt_513/ptr_deref_500_Update/word_access_complete/word_0/cr
      -- CP-element group 231: 	 branch_block_stmt_239/merge_stmt_350_PhiAck/$exit
      -- CP-element group 231: 	 branch_block_stmt_239/merge_stmt_350_PhiAck/phi_stmt_351_ack
      -- 
    phi_stmt_351_ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_351_ack_0, ack => zeropad3D_CP_676_elements(231)); -- 
    req_974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => array_obj_ref_363_index_offset_req_0); -- 
    req_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => array_obj_ref_363_index_offset_req_1); -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => addr_of_364_final_reg_req_1); -- 
    rr_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => RPIPE_zeropad_input_pipe_367_inst_req_0); -- 
    cr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_371_inst_req_1); -- 
    cr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_384_inst_req_1); -- 
    cr_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_402_inst_req_1); -- 
    cr_1106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_420_inst_req_1); -- 
    cr_1134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_438_inst_req_1); -- 
    cr_1162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_456_inst_req_1); -- 
    cr_1190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_474_inst_req_1); -- 
    cr_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => type_cast_492_inst_req_1); -- 
    cr_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(231), ack => ptr_deref_500_store_0_req_1); -- 
    -- CP-element group 232:  merge  fork  transition  place  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	26 
    -- CP-element group 232: 	75 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	77 
    -- CP-element group 232: 	78 
    -- CP-element group 232: 	80 
    -- CP-element group 232: 	81 
    -- CP-element group 232: 	95 
    -- CP-element group 232: 	109 
    -- CP-element group 232: 	123 
    -- CP-element group 232: 	137 
    -- CP-element group 232: 	151 
    -- CP-element group 232: 	165 
    -- CP-element group 232: 	179 
    -- CP-element group 232:  members (40) 
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699__entry__
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/merge_stmt_522__exit__
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block2_starting_574_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block3_starting_595_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block4_starting_616_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block5_starting_637_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_update_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Sample/crr
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Update/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/call_stmt_525_Update/ccr
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_update_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Update/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/type_cast_530_Update/cr
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block0_starting_532_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block1_starting_553_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block6_starting_658_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_239/call_stmt_525_to_assign_stmt_699/WPIPE_Block7_starting_679_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_239/merge_stmt_522_PhiAck/dummy
      -- CP-element group 232: 	 branch_block_stmt_239/merge_stmt_522_PhiAck/$exit
      -- CP-element group 232: 	 branch_block_stmt_239/merge_stmt_522_PhiReqMerge
      -- CP-element group 232: 	 branch_block_stmt_239/merge_stmt_522_PhiAck/$entry
      -- 
    req_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block3_starting_595_inst_req_0); -- 
    req_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block2_starting_574_inst_req_0); -- 
    req_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block4_starting_616_inst_req_0); -- 
    req_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block5_starting_637_inst_req_0); -- 
    crr_1299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => call_stmt_525_call_req_0); -- 
    ccr_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => call_stmt_525_call_req_1); -- 
    cr_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => type_cast_530_inst_req_1); -- 
    req_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block0_starting_532_inst_req_0); -- 
    req_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block1_starting_553_inst_req_0); -- 
    req_1915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block6_starting_658_inst_req_0); -- 
    req_2013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => WPIPE_Block7_starting_679_inst_req_0); -- 
    zeropad3D_CP_676_elements(232) <= OrReduce(zeropad3D_CP_676_elements(26) & zeropad3D_CP_676_elements(75));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_362_resized : std_logic_vector(13 downto 0);
    signal R_indvar_362_scaled : std_logic_vector(13 downto 0);
    signal add31_408 : std_logic_vector(63 downto 0);
    signal add37_426 : std_logic_vector(63 downto 0);
    signal add43_444 : std_logic_vector(63 downto 0);
    signal add49_462 : std_logic_vector(63 downto 0);
    signal add55_480 : std_logic_vector(63 downto 0);
    signal add61_498 : std_logic_vector(63 downto 0);
    signal add_390 : std_logic_vector(63 downto 0);
    signal array_obj_ref_363_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_363_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_365 : std_logic_vector(31 downto 0);
    signal call125_703 : std_logic_vector(7 downto 0);
    signal call128_706 : std_logic_vector(7 downto 0);
    signal call131_709 : std_logic_vector(7 downto 0);
    signal call134_712 : std_logic_vector(7 downto 0);
    signal call137_715 : std_logic_vector(7 downto 0);
    signal call140_718 : std_logic_vector(7 downto 0);
    signal call143_721 : std_logic_vector(7 downto 0);
    signal call146_724 : std_logic_vector(7 downto 0);
    signal call149_727 : std_logic_vector(63 downto 0);
    signal call1_245 : std_logic_vector(7 downto 0);
    signal call20_368 : std_logic_vector(7 downto 0);
    signal call23_381 : std_logic_vector(7 downto 0);
    signal call28_399 : std_logic_vector(7 downto 0);
    signal call2_248 : std_logic_vector(7 downto 0);
    signal call34_417 : std_logic_vector(7 downto 0);
    signal call3_251 : std_logic_vector(7 downto 0);
    signal call40_435 : std_logic_vector(7 downto 0);
    signal call46_453 : std_logic_vector(7 downto 0);
    signal call4_254 : std_logic_vector(7 downto 0);
    signal call52_471 : std_logic_vector(7 downto 0);
    signal call58_489 : std_logic_vector(7 downto 0);
    signal call5_257 : std_logic_vector(7 downto 0);
    signal call66_525 : std_logic_vector(63 downto 0);
    signal call6_260 : std_logic_vector(7 downto 0);
    signal call7_263 : std_logic_vector(7 downto 0);
    signal call8_266 : std_logic_vector(7 downto 0);
    signal call_242 : std_logic_vector(7 downto 0);
    signal cmp166_300 : std_logic_vector(0 downto 0);
    signal conv10_274 : std_logic_vector(63 downto 0);
    signal conv12_278 : std_logic_vector(63 downto 0);
    signal conv150_732 : std_logic_vector(63 downto 0);
    signal conv156_745 : std_logic_vector(31 downto 0);
    signal conv158_749 : std_logic_vector(31 downto 0);
    signal conv161_753 : std_logic_vector(31 downto 0);
    signal conv21_372 : std_logic_vector(63 downto 0);
    signal conv25_385 : std_logic_vector(63 downto 0);
    signal conv30_403 : std_logic_vector(63 downto 0);
    signal conv36_421 : std_logic_vector(63 downto 0);
    signal conv42_439 : std_logic_vector(63 downto 0);
    signal conv48_457 : std_logic_vector(63 downto 0);
    signal conv54_475 : std_logic_vector(63 downto 0);
    signal conv60_493 : std_logic_vector(63 downto 0);
    signal conv67_531 : std_logic_vector(63 downto 0);
    signal conv_270 : std_logic_vector(63 downto 0);
    signal exitcond8_513 : std_logic_vector(0 downto 0);
    signal indvar_351 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_508 : std_logic_vector(63 downto 0);
    signal mul13_288 : std_logic_vector(63 downto 0);
    signal mul159_758 : std_logic_vector(31 downto 0);
    signal mul162_763 : std_logic_vector(31 downto 0);
    signal mul_283 : std_logic_vector(63 downto 0);
    signal ptr_deref_500_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_500_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_500_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_500_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_500_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_500_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl27_396 : std_logic_vector(63 downto 0);
    signal shl33_414 : std_logic_vector(63 downto 0);
    signal shl39_432 : std_logic_vector(63 downto 0);
    signal shl45_450 : std_logic_vector(63 downto 0);
    signal shl51_468 : std_logic_vector(63 downto 0);
    signal shl57_486 : std_logic_vector(63 downto 0);
    signal shl_378 : std_logic_vector(63 downto 0);
    signal shr165x_xmask_294 : std_logic_vector(63 downto 0);
    signal sub_737 : std_logic_vector(63 downto 0);
    signal tmp1_315 : std_logic_vector(63 downto 0);
    signal tmp2_320 : std_logic_vector(63 downto 0);
    signal tmp3_324 : std_logic_vector(63 downto 0);
    signal tmp4_329 : std_logic_vector(63 downto 0);
    signal tmp5_335 : std_logic_vector(63 downto 0);
    signal tmp6_341 : std_logic_vector(0 downto 0);
    signal tmp_311 : std_logic_vector(63 downto 0);
    signal type_cast_292_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_298_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_333_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_339_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_355_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_357_wire : std_logic_vector(63 downto 0);
    signal type_cast_376_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_412_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_430_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_466_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_484_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_506_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_529_wire : std_logic_vector(63 downto 0);
    signal type_cast_730_wire : std_logic_vector(63 downto 0);
    signal umax7_348 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_363_constant_part_of_offset <= "00000000000000";
    array_obj_ref_363_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_363_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_363_resized_base_address <= "00000000000000";
    ptr_deref_500_word_offset_0 <= "00000000000000";
    type_cast_292_wire_constant <= "0000000000000000000000000000000000000000111111111111111111111100";
    type_cast_298_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_339_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_355_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_376_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_412_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_430_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_448_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_466_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_484_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_506_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_351: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_355_wire_constant & type_cast_357_wire;
      req <= phi_stmt_351_req_0 & phi_stmt_351_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_351",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_351_ack_0,
          idata => idata,
          odata => indvar_351,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_351
    -- flow-through select operator MUX_347_inst
    umax7_348 <= tmp5_335 when (tmp6_341(0) /=  '0') else type_cast_346_wire_constant;
    addr_of_364_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_364_final_reg_req_0;
      addr_of_364_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_364_final_reg_req_1;
      addr_of_364_final_reg_ack_1<= rack(0);
      addr_of_364_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_364_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_363_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_273_inst_req_0;
      type_cast_273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_273_inst_req_1;
      type_cast_273_inst_ack_1<= rack(0);
      type_cast_273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_277_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_277_inst_req_0;
      type_cast_277_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_277_inst_req_1;
      type_cast_277_inst_ack_1<= rack(0);
      type_cast_277_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_277_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_310_inst_req_0;
      type_cast_310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_310_inst_req_1;
      type_cast_310_inst_ack_1<= rack(0);
      type_cast_310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_314_inst_req_0;
      type_cast_314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_314_inst_req_1;
      type_cast_314_inst_ack_1<= rack(0);
      type_cast_314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_323_inst_req_0;
      type_cast_323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_323_inst_req_1;
      type_cast_323_inst_ack_1<= rack(0);
      type_cast_323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_324,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_508,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_357_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_384_inst_req_0;
      type_cast_384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_384_inst_req_1;
      type_cast_384_inst_ack_1<= rack(0);
      type_cast_384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv25_385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_402_inst_req_0;
      type_cast_402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_402_inst_req_1;
      type_cast_402_inst_ack_1<= rack(0);
      type_cast_402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_420_inst_req_0;
      type_cast_420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_420_inst_req_1;
      type_cast_420_inst_ack_1<= rack(0);
      type_cast_420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call34_417,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_438_inst_req_0;
      type_cast_438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_438_inst_req_1;
      type_cast_438_inst_ack_1<= rack(0);
      type_cast_438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_456_inst_req_0;
      type_cast_456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_456_inst_req_1;
      type_cast_456_inst_ack_1<= rack(0);
      type_cast_456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_474_inst_req_0;
      type_cast_474_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_474_inst_req_1;
      type_cast_474_inst_ack_1<= rack(0);
      type_cast_474_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_474_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call52_471,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_492_inst_req_0;
      type_cast_492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_492_inst_req_1;
      type_cast_492_inst_ack_1<= rack(0);
      type_cast_492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call58_489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_530_inst_req_0;
      type_cast_530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_530_inst_req_1;
      type_cast_530_inst_ack_1<= rack(0);
      type_cast_530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_529_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_531,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_730_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_744_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_744_inst_req_0;
      type_cast_744_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_744_inst_req_1;
      type_cast_744_inst_ack_1<= rack(0);
      type_cast_744_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_744_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv156_745,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_748_inst_req_0;
      type_cast_748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_748_inst_req_1;
      type_cast_748_inst_ack_1<= rack(0);
      type_cast_748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_752_inst_req_0;
      type_cast_752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_752_inst_req_1;
      type_cast_752_inst_ack_1<= rack(0);
      type_cast_752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call8_266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_753,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_363_index_1_rename
    process(R_indvar_362_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_362_resized;
      ov(13 downto 0) := iv;
      R_indvar_362_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_index_1_resize
    process(indvar_351) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_351;
      ov := iv(13 downto 0);
      R_indvar_362_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_root_address_inst
    process(array_obj_ref_363_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_363_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_363_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_addr_0
    process(ptr_deref_500_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_500_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_base_resize
    process(arrayidx_365) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_365;
      ov := iv(13 downto 0);
      ptr_deref_500_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_gather_scatter
    process(add61_498) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add61_498;
      ov(63 downto 0) := iv;
      ptr_deref_500_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_root_address_inst
    process(ptr_deref_500_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_500_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_301_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp166_300;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_301_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_301_branch_req_0,
          ack0 => if_stmt_301_branch_ack_0,
          ack1 => if_stmt_301_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_514_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond8_513;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_514_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_514_branch_req_0,
          ack0 => if_stmt_514_branch_ack_0,
          ack1 => if_stmt_514_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_507_inst
    process(indvar_351) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_351, type_cast_506_wire_constant, tmp_var);
      indvarx_xnext_508 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_293_inst
    process(mul13_288) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul13_288, type_cast_292_wire_constant, tmp_var);
      shr165x_xmask_294 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_299_inst
    process(shr165x_xmask_294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr165x_xmask_294, type_cast_298_wire_constant, tmp_var);
      cmp166_300 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_512_inst
    process(indvarx_xnext_508, umax7_348) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_508, umax7_348, tmp_var);
      exitcond8_513 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_334_inst
    process(tmp4_329) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_329, type_cast_333_wire_constant, tmp_var);
      tmp5_335 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_757_inst
    process(conv158_749, conv156_745) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv158_749, conv156_745, tmp_var);
      mul159_758 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_762_inst
    process(mul159_758, conv161_753) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul159_758, conv161_753, tmp_var);
      mul162_763 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_282_inst
    process(conv10_274, conv_270) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv10_274, conv_270, tmp_var);
      mul_283 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_287_inst
    process(mul_283, conv12_278) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_283, conv12_278, tmp_var);
      mul13_288 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_319_inst
    process(tmp_311, tmp1_315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_311, tmp1_315, tmp_var);
      tmp2_320 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_328_inst
    process(tmp2_320, tmp3_324) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_320, tmp3_324, tmp_var);
      tmp4_329 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_389_inst
    process(shl_378, conv25_385) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_378, conv25_385, tmp_var);
      add_390 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_407_inst
    process(shl27_396, conv30_403) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_396, conv30_403, tmp_var);
      add31_408 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_425_inst
    process(shl33_414, conv36_421) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl33_414, conv36_421, tmp_var);
      add37_426 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_443_inst
    process(shl39_432, conv42_439) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl39_432, conv42_439, tmp_var);
      add43_444 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_461_inst
    process(shl45_450, conv48_457) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_450, conv48_457, tmp_var);
      add49_462 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_479_inst
    process(shl51_468, conv54_475) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl51_468, conv54_475, tmp_var);
      add55_480 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_497_inst
    process(shl57_486, conv60_493) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl57_486, conv60_493, tmp_var);
      add61_498 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_377_inst
    process(conv21_372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv21_372, type_cast_376_wire_constant, tmp_var);
      shl_378 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_395_inst
    process(add_390) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_390, type_cast_394_wire_constant, tmp_var);
      shl27_396 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_413_inst
    process(add31_408) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add31_408, type_cast_412_wire_constant, tmp_var);
      shl33_414 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_431_inst
    process(add37_426) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add37_426, type_cast_430_wire_constant, tmp_var);
      shl39_432 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_449_inst
    process(add43_444) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add43_444, type_cast_448_wire_constant, tmp_var);
      shl45_450 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_467_inst
    process(add49_462) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add49_462, type_cast_466_wire_constant, tmp_var);
      shl51_468 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_485_inst
    process(add55_480) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add55_480, type_cast_484_wire_constant, tmp_var);
      shl57_486 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_736_inst
    process(conv150_732, conv67_531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv150_732, conv67_531, tmp_var);
      sub_737 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_340_inst
    process(tmp5_335) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp5_335, type_cast_339_wire_constant, tmp_var);
      tmp6_341 <= tmp_var; --
    end process;
    -- shared split operator group (27) : array_obj_ref_363_index_offset 
    ApIntAdd_group_27: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_362_scaled;
      array_obj_ref_363_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_363_index_offset_req_0;
      array_obj_ref_363_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_363_index_offset_req_1;
      array_obj_ref_363_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_27_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- unary operator type_cast_529_inst
    process(call66_525) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call66_525, tmp_var);
      type_cast_529_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_730_inst
    process(call149_727) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call149_727, tmp_var);
      type_cast_730_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_500_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_500_store_0_req_0;
      ptr_deref_500_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_500_store_0_req_1;
      ptr_deref_500_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_500_word_address_0;
      data_in <= ptr_deref_500_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_complete_702_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_complete_702_inst_req_0;
      RPIPE_Block0_complete_702_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_complete_702_inst_req_1;
      RPIPE_Block0_complete_702_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call125_703 <= data_out(7 downto 0);
      Block0_complete_read_0_gI: SplitGuardInterface generic map(name => "Block0_complete_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_complete_read_0: InputPortRevised -- 
        generic map ( name => "Block0_complete_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_complete_pipe_read_req(0),
          oack => Block0_complete_pipe_read_ack(0),
          odata => Block0_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_complete_705_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_complete_705_inst_req_0;
      RPIPE_Block1_complete_705_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_complete_705_inst_req_1;
      RPIPE_Block1_complete_705_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call128_706 <= data_out(7 downto 0);
      Block1_complete_read_1_gI: SplitGuardInterface generic map(name => "Block1_complete_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_complete_read_1: InputPortRevised -- 
        generic map ( name => "Block1_complete_read_1", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_complete_pipe_read_req(0),
          oack => Block1_complete_pipe_read_ack(0),
          odata => Block1_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_complete_708_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_complete_708_inst_req_0;
      RPIPE_Block2_complete_708_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_complete_708_inst_req_1;
      RPIPE_Block2_complete_708_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call131_709 <= data_out(7 downto 0);
      Block2_complete_read_2_gI: SplitGuardInterface generic map(name => "Block2_complete_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_complete_read_2: InputPortRevised -- 
        generic map ( name => "Block2_complete_read_2", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_complete_pipe_read_req(0),
          oack => Block2_complete_pipe_read_ack(0),
          odata => Block2_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_complete_711_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_complete_711_inst_req_0;
      RPIPE_Block3_complete_711_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_complete_711_inst_req_1;
      RPIPE_Block3_complete_711_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call134_712 <= data_out(7 downto 0);
      Block3_complete_read_3_gI: SplitGuardInterface generic map(name => "Block3_complete_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_complete_read_3: InputPortRevised -- 
        generic map ( name => "Block3_complete_read_3", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_complete_pipe_read_req(0),
          oack => Block3_complete_pipe_read_ack(0),
          odata => Block3_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_Block4_complete_714_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block4_complete_714_inst_req_0;
      RPIPE_Block4_complete_714_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block4_complete_714_inst_req_1;
      RPIPE_Block4_complete_714_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call137_715 <= data_out(7 downto 0);
      Block4_complete_read_4_gI: SplitGuardInterface generic map(name => "Block4_complete_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block4_complete_read_4: InputPortRevised -- 
        generic map ( name => "Block4_complete_read_4", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block4_complete_pipe_read_req(0),
          oack => Block4_complete_pipe_read_ack(0),
          odata => Block4_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_Block5_complete_717_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block5_complete_717_inst_req_0;
      RPIPE_Block5_complete_717_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block5_complete_717_inst_req_1;
      RPIPE_Block5_complete_717_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call140_718 <= data_out(7 downto 0);
      Block5_complete_read_5_gI: SplitGuardInterface generic map(name => "Block5_complete_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block5_complete_read_5: InputPortRevised -- 
        generic map ( name => "Block5_complete_read_5", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block5_complete_pipe_read_req(0),
          oack => Block5_complete_pipe_read_ack(0),
          odata => Block5_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_Block6_complete_720_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block6_complete_720_inst_req_0;
      RPIPE_Block6_complete_720_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block6_complete_720_inst_req_1;
      RPIPE_Block6_complete_720_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call143_721 <= data_out(7 downto 0);
      Block6_complete_read_6_gI: SplitGuardInterface generic map(name => "Block6_complete_read_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block6_complete_read_6: InputPortRevised -- 
        generic map ( name => "Block6_complete_read_6", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block6_complete_pipe_read_req(0),
          oack => Block6_complete_pipe_read_ack(0),
          odata => Block6_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_Block7_complete_723_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block7_complete_723_inst_req_0;
      RPIPE_Block7_complete_723_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block7_complete_723_inst_req_1;
      RPIPE_Block7_complete_723_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call146_724 <= data_out(7 downto 0);
      Block7_complete_read_7_gI: SplitGuardInterface generic map(name => "Block7_complete_read_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block7_complete_read_7: InputPortRevised -- 
        generic map ( name => "Block7_complete_read_7", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block7_complete_pipe_read_req(0),
          oack => Block7_complete_pipe_read_ack(0),
          odata => Block7_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_zeropad_input_pipe_470_inst RPIPE_zeropad_input_pipe_398_inst RPIPE_zeropad_input_pipe_452_inst RPIPE_zeropad_input_pipe_380_inst RPIPE_zeropad_input_pipe_434_inst RPIPE_zeropad_input_pipe_265_inst RPIPE_zeropad_input_pipe_262_inst RPIPE_zeropad_input_pipe_259_inst RPIPE_zeropad_input_pipe_488_inst RPIPE_zeropad_input_pipe_256_inst RPIPE_zeropad_input_pipe_253_inst RPIPE_zeropad_input_pipe_367_inst RPIPE_zeropad_input_pipe_250_inst RPIPE_zeropad_input_pipe_416_inst RPIPE_zeropad_input_pipe_247_inst RPIPE_zeropad_input_pipe_244_inst RPIPE_zeropad_input_pipe_241_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(135 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 16 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_470_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_398_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_452_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_380_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_434_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_265_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_262_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_259_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_488_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_256_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_253_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_367_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_250_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_416_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_247_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_244_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_241_inst_req_0;
      RPIPE_zeropad_input_pipe_470_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_398_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_452_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_380_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_434_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_265_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_262_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_259_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_488_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_256_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_253_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_367_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_250_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_416_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_247_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_244_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_241_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_470_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_398_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_452_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_380_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_434_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_265_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_262_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_259_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_488_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_256_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_253_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_367_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_250_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_416_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_247_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_244_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_241_inst_req_1;
      RPIPE_zeropad_input_pipe_470_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_398_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_452_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_380_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_434_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_265_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_262_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_259_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_488_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_256_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_253_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_367_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_250_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_416_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_247_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_244_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_241_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      call52_471 <= data_out(135 downto 128);
      call28_399 <= data_out(127 downto 120);
      call46_453 <= data_out(119 downto 112);
      call23_381 <= data_out(111 downto 104);
      call40_435 <= data_out(103 downto 96);
      call8_266 <= data_out(95 downto 88);
      call7_263 <= data_out(87 downto 80);
      call6_260 <= data_out(79 downto 72);
      call58_489 <= data_out(71 downto 64);
      call5_257 <= data_out(63 downto 56);
      call4_254 <= data_out(55 downto 48);
      call20_368 <= data_out(47 downto 40);
      call3_251 <= data_out(39 downto 32);
      call34_417 <= data_out(31 downto 24);
      call2_248 <= data_out(23 downto 16);
      call1_245 <= data_out(15 downto 8);
      call_242 <= data_out(7 downto 0);
      zeropad_input_pipe_read_8_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_8_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_8: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_8", data_width => 8,  num_reqs => 17,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared outport operator group (0) : WPIPE_Block0_starting_547_inst WPIPE_Block0_starting_550_inst WPIPE_Block0_starting_544_inst WPIPE_Block0_starting_541_inst WPIPE_Block0_starting_532_inst WPIPE_Block0_starting_538_inst WPIPE_Block0_starting_535_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block0_starting_547_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_starting_550_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_starting_544_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_starting_541_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_starting_532_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_starting_538_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_starting_535_inst_req_0;
      WPIPE_Block0_starting_547_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_starting_550_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_starting_544_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_starting_541_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_starting_532_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_starting_538_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_starting_535_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block0_starting_547_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_starting_550_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_starting_544_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_starting_541_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_starting_532_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_starting_538_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_starting_535_inst_req_1;
      WPIPE_Block0_starting_547_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_starting_550_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_starting_544_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_starting_541_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_starting_532_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_starting_538_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_starting_535_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call8_266 & call5_257 & call7_263 & call6_260 & call2_248 & call4_254 & call3_251;
      Block0_starting_write_0_gI: SplitGuardInterface generic map(name => "Block0_starting_write_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_starting_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_starting_pipe_write_req(0),
          oack => Block0_starting_pipe_write_ack(0),
          odata => Block0_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_starting_571_inst WPIPE_Block1_starting_568_inst WPIPE_Block1_starting_565_inst WPIPE_Block1_starting_562_inst WPIPE_Block1_starting_559_inst WPIPE_Block1_starting_556_inst WPIPE_Block1_starting_553_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block1_starting_571_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_starting_568_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_starting_565_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_starting_562_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_starting_559_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_starting_556_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_starting_553_inst_req_0;
      WPIPE_Block1_starting_571_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_starting_568_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_starting_565_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_starting_562_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_starting_559_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_starting_556_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_starting_553_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block1_starting_571_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_starting_568_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_starting_565_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_starting_562_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_starting_559_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_starting_556_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_starting_553_inst_req_1;
      WPIPE_Block1_starting_571_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_starting_568_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_starting_565_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_starting_562_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_starting_559_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_starting_556_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_starting_553_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call5_257 & call8_266 & call7_263 & call6_260 & call4_254 & call3_251 & call2_248;
      Block1_starting_write_1_gI: SplitGuardInterface generic map(name => "Block1_starting_write_1_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_starting_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_starting_pipe_write_req(0),
          oack => Block1_starting_pipe_write_ack(0),
          odata => Block1_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_starting_592_inst WPIPE_Block2_starting_589_inst WPIPE_Block2_starting_586_inst WPIPE_Block2_starting_583_inst WPIPE_Block2_starting_580_inst WPIPE_Block2_starting_577_inst WPIPE_Block2_starting_574_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block2_starting_592_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_starting_589_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_starting_586_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_starting_583_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_starting_580_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_starting_577_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_starting_574_inst_req_0;
      WPIPE_Block2_starting_592_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_starting_589_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_starting_586_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_starting_583_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_starting_580_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_starting_577_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_starting_574_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block2_starting_592_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_starting_589_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_starting_586_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_starting_583_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_starting_580_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_starting_577_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_starting_574_inst_req_1;
      WPIPE_Block2_starting_592_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_starting_589_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_starting_586_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_starting_583_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_starting_580_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_starting_577_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_starting_574_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call5_257 & call8_266 & call7_263 & call6_260 & call4_254 & call3_251 & call2_248;
      Block2_starting_write_2_gI: SplitGuardInterface generic map(name => "Block2_starting_write_2_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_starting_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_starting_pipe_write_req(0),
          oack => Block2_starting_pipe_write_ack(0),
          odata => Block2_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_starting_595_inst WPIPE_Block3_starting_598_inst WPIPE_Block3_starting_601_inst WPIPE_Block3_starting_604_inst WPIPE_Block3_starting_607_inst WPIPE_Block3_starting_613_inst WPIPE_Block3_starting_610_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block3_starting_595_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_starting_598_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_starting_601_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_starting_604_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_starting_607_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_starting_613_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_starting_610_inst_req_0;
      WPIPE_Block3_starting_595_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_starting_598_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_starting_601_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_starting_604_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_starting_607_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_starting_613_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_starting_610_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block3_starting_595_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_starting_598_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_starting_601_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_starting_604_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_starting_607_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_starting_613_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_starting_610_inst_req_1;
      WPIPE_Block3_starting_595_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_starting_598_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_starting_601_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_starting_604_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_starting_607_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_starting_613_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_starting_610_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call2_248 & call3_251 & call4_254 & call6_260 & call7_263 & call5_257 & call8_266;
      Block3_starting_write_3_gI: SplitGuardInterface generic map(name => "Block3_starting_write_3_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_starting_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_starting_pipe_write_req(0),
          oack => Block3_starting_pipe_write_ack(0),
          odata => Block3_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_Block4_starting_619_inst WPIPE_Block4_starting_622_inst WPIPE_Block4_starting_634_inst WPIPE_Block4_starting_631_inst WPIPE_Block4_starting_628_inst WPIPE_Block4_starting_625_inst WPIPE_Block4_starting_616_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block4_starting_619_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block4_starting_622_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block4_starting_634_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block4_starting_631_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block4_starting_628_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block4_starting_625_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block4_starting_616_inst_req_0;
      WPIPE_Block4_starting_619_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block4_starting_622_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block4_starting_634_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block4_starting_631_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block4_starting_628_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block4_starting_625_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block4_starting_616_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block4_starting_619_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block4_starting_622_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block4_starting_634_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block4_starting_631_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block4_starting_628_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block4_starting_625_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block4_starting_616_inst_req_1;
      WPIPE_Block4_starting_619_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block4_starting_622_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block4_starting_634_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block4_starting_631_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block4_starting_628_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block4_starting_625_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block4_starting_616_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call3_251 & call4_254 & call5_257 & call8_266 & call7_263 & call6_260 & call2_248;
      Block4_starting_write_4_gI: SplitGuardInterface generic map(name => "Block4_starting_write_4_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block4_starting_write_4: OutputPortRevised -- 
        generic map ( name => "Block4_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block4_starting_pipe_write_req(0),
          oack => Block4_starting_pipe_write_ack(0),
          odata => Block4_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_Block5_starting_655_inst WPIPE_Block5_starting_652_inst WPIPE_Block5_starting_649_inst WPIPE_Block5_starting_646_inst WPIPE_Block5_starting_643_inst WPIPE_Block5_starting_640_inst WPIPE_Block5_starting_637_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block5_starting_655_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block5_starting_652_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block5_starting_649_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block5_starting_646_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block5_starting_643_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block5_starting_640_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block5_starting_637_inst_req_0;
      WPIPE_Block5_starting_655_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block5_starting_652_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block5_starting_649_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block5_starting_646_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block5_starting_643_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block5_starting_640_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block5_starting_637_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block5_starting_655_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block5_starting_652_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block5_starting_649_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block5_starting_646_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block5_starting_643_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block5_starting_640_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block5_starting_637_inst_req_1;
      WPIPE_Block5_starting_655_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block5_starting_652_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block5_starting_649_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block5_starting_646_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block5_starting_643_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block5_starting_640_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block5_starting_637_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call5_257 & call8_266 & call7_263 & call6_260 & call4_254 & call3_251 & call2_248;
      Block5_starting_write_5_gI: SplitGuardInterface generic map(name => "Block5_starting_write_5_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block5_starting_write_5: OutputPortRevised -- 
        generic map ( name => "Block5_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block5_starting_pipe_write_req(0),
          oack => Block5_starting_pipe_write_ack(0),
          odata => Block5_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_Block6_starting_676_inst WPIPE_Block6_starting_673_inst WPIPE_Block6_starting_670_inst WPIPE_Block6_starting_667_inst WPIPE_Block6_starting_664_inst WPIPE_Block6_starting_661_inst WPIPE_Block6_starting_658_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block6_starting_676_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block6_starting_673_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block6_starting_670_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block6_starting_667_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block6_starting_664_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block6_starting_661_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block6_starting_658_inst_req_0;
      WPIPE_Block6_starting_676_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block6_starting_673_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block6_starting_670_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block6_starting_667_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block6_starting_664_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block6_starting_661_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block6_starting_658_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block6_starting_676_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block6_starting_673_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block6_starting_670_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block6_starting_667_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block6_starting_664_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block6_starting_661_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block6_starting_658_inst_req_1;
      WPIPE_Block6_starting_676_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block6_starting_673_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block6_starting_670_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block6_starting_667_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block6_starting_664_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block6_starting_661_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block6_starting_658_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call5_257 & call8_266 & call7_263 & call6_260 & call4_254 & call3_251 & call2_248;
      Block6_starting_write_6_gI: SplitGuardInterface generic map(name => "Block6_starting_write_6_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block6_starting_write_6: OutputPortRevised -- 
        generic map ( name => "Block6_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block6_starting_pipe_write_req(0),
          oack => Block6_starting_pipe_write_ack(0),
          odata => Block6_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_Block7_starting_685_inst WPIPE_Block7_starting_682_inst WPIPE_Block7_starting_679_inst WPIPE_Block7_starting_697_inst WPIPE_Block7_starting_694_inst WPIPE_Block7_starting_691_inst WPIPE_Block7_starting_688_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block7_starting_685_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block7_starting_682_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block7_starting_679_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block7_starting_697_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block7_starting_694_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block7_starting_691_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block7_starting_688_inst_req_0;
      WPIPE_Block7_starting_685_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block7_starting_682_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block7_starting_679_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block7_starting_697_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block7_starting_694_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block7_starting_691_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block7_starting_688_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block7_starting_685_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block7_starting_682_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block7_starting_679_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block7_starting_697_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block7_starting_694_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block7_starting_691_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block7_starting_688_inst_req_1;
      WPIPE_Block7_starting_685_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block7_starting_682_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block7_starting_679_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block7_starting_697_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block7_starting_694_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block7_starting_691_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block7_starting_688_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call4_254 & call3_251 & call2_248 & call5_257 & call8_266 & call7_263 & call6_260;
      Block7_starting_write_7_gI: SplitGuardInterface generic map(name => "Block7_starting_write_7_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block7_starting_write_7: OutputPortRevised -- 
        generic map ( name => "Block7_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block7_starting_pipe_write_req(0),
          oack => Block7_starting_pipe_write_ack(0),
          odata => Block7_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- shared outport operator group (8) : WPIPE_elapsed_time_pipe_738_inst 
    OutportGroup_8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_738_inst_req_0;
      WPIPE_elapsed_time_pipe_738_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_738_inst_req_1;
      WPIPE_elapsed_time_pipe_738_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_737;
      elapsed_time_pipe_write_8_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_8: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- shared call operator group (0) : call_stmt_525_call call_stmt_727_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_525_call_req_0;
      reqL_unguarded(0) <= call_stmt_727_call_req_0;
      call_stmt_525_call_ack_0 <= ackL_unguarded(1);
      call_stmt_727_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_525_call_req_1;
      reqR_unguarded(0) <= call_stmt_727_call_req_1;
      call_stmt_525_call_ack_1 <= ackR_unguarded(1);
      call_stmt_727_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call66_525 <= data_out(127 downto 64);
      call149_727 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_765_call 
    sendOutput_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_765_call_req_0;
      call_stmt_765_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_765_call_req_1;
      call_stmt_765_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul162_763;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          dataR => sendOutput_call_data(31 downto 0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_A is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_A;
architecture zeropad3D_A_arch of zeropad3D_A is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_A_CP_2408_start: Boolean;
  signal zeropad3D_A_CP_2408_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_starting_776_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_776_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_779_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_776_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal phi_stmt_910_req_1 : boolean;
  signal RPIPE_Block0_starting_779_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_779_inst_ack_0 : boolean;
  signal if_stmt_1239_branch_ack_0 : boolean;
  signal if_stmt_1182_branch_ack_1 : boolean;
  signal type_cast_1206_inst_ack_0 : boolean;
  signal if_stmt_1182_branch_req_0 : boolean;
  signal if_stmt_1239_branch_ack_1 : boolean;
  signal RPIPE_Block0_starting_773_inst_req_0 : boolean;
  signal type_cast_1206_inst_req_0 : boolean;
  signal type_cast_1149_inst_ack_1 : boolean;
  signal type_cast_1149_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_773_inst_ack_0 : boolean;
  signal addr_of_1156_final_reg_ack_1 : boolean;
  signal RPIPE_Block0_starting_773_inst_req_1 : boolean;
  signal type_cast_909_inst_req_0 : boolean;
  signal type_cast_909_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_773_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_779_inst_ack_1 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal array_obj_ref_1155_index_offset_req_0 : boolean;
  signal RPIPE_Block0_starting_776_inst_req_1 : boolean;
  signal type_cast_1149_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_782_inst_req_0 : boolean;
  signal type_cast_1256_inst_ack_1 : boolean;
  signal if_stmt_1182_branch_ack_0 : boolean;
  signal type_cast_1249_inst_ack_1 : boolean;
  signal phi_stmt_1253_req_1 : boolean;
  signal type_cast_1256_inst_req_1 : boolean;
  signal type_cast_1249_inst_ack_0 : boolean;
  signal type_cast_1249_inst_req_0 : boolean;
  signal array_obj_ref_1155_index_offset_ack_0 : boolean;
  signal type_cast_1262_inst_ack_0 : boolean;
  signal type_cast_1262_inst_req_0 : boolean;
  signal type_cast_1264_inst_req_0 : boolean;
  signal type_cast_1206_inst_req_1 : boolean;
  signal type_cast_1264_inst_ack_0 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal type_cast_1206_inst_ack_1 : boolean;
  signal array_obj_ref_1155_index_offset_req_1 : boolean;
  signal array_obj_ref_1155_index_offset_ack_1 : boolean;
  signal type_cast_1264_inst_req_1 : boolean;
  signal WPIPE_Block0_complete_1269_inst_req_0 : boolean;
  signal type_cast_1264_inst_ack_1 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal phi_stmt_1253_req_0 : boolean;
  signal WPIPE_Block0_complete_1269_inst_ack_0 : boolean;
  signal type_cast_1262_inst_req_1 : boolean;
  signal type_cast_1262_inst_ack_1 : boolean;
  signal phi_stmt_1259_req_0 : boolean;
  signal WPIPE_Block0_complete_1269_inst_req_1 : boolean;
  signal type_cast_1249_inst_req_1 : boolean;
  signal WPIPE_Block0_complete_1269_inst_ack_1 : boolean;
  signal phi_stmt_1259_req_1 : boolean;
  signal phi_stmt_1246_req_0 : boolean;
  signal type_cast_1215_inst_req_0 : boolean;
  signal type_cast_1256_inst_req_0 : boolean;
  signal type_cast_1258_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_782_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_782_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_782_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_785_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_785_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_785_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_785_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_788_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_788_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_788_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_788_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_791_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_791_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_791_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_791_inst_ack_1 : boolean;
  signal type_cast_796_inst_req_0 : boolean;
  signal type_cast_796_inst_ack_0 : boolean;
  signal type_cast_796_inst_req_1 : boolean;
  signal type_cast_796_inst_ack_1 : boolean;
  signal type_cast_800_inst_req_0 : boolean;
  signal type_cast_800_inst_ack_0 : boolean;
  signal type_cast_800_inst_req_1 : boolean;
  signal type_cast_800_inst_ack_1 : boolean;
  signal type_cast_804_inst_req_0 : boolean;
  signal type_cast_804_inst_ack_0 : boolean;
  signal type_cast_804_inst_req_1 : boolean;
  signal type_cast_804_inst_ack_1 : boolean;
  signal type_cast_808_inst_req_0 : boolean;
  signal type_cast_808_inst_ack_0 : boolean;
  signal type_cast_808_inst_req_1 : boolean;
  signal type_cast_808_inst_ack_1 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal type_cast_821_inst_req_0 : boolean;
  signal type_cast_821_inst_ack_0 : boolean;
  signal type_cast_821_inst_req_1 : boolean;
  signal type_cast_821_inst_ack_1 : boolean;
  signal type_cast_857_inst_req_0 : boolean;
  signal type_cast_857_inst_ack_0 : boolean;
  signal type_cast_857_inst_req_1 : boolean;
  signal type_cast_857_inst_ack_1 : boolean;
  signal type_cast_928_inst_req_0 : boolean;
  signal type_cast_928_inst_ack_0 : boolean;
  signal type_cast_928_inst_req_1 : boolean;
  signal type_cast_928_inst_ack_1 : boolean;
  signal if_stmt_955_branch_req_0 : boolean;
  signal if_stmt_955_branch_ack_1 : boolean;
  signal if_stmt_955_branch_ack_0 : boolean;
  signal type_cast_965_inst_req_0 : boolean;
  signal type_cast_965_inst_ack_0 : boolean;
  signal type_cast_965_inst_req_1 : boolean;
  signal type_cast_965_inst_ack_1 : boolean;
  signal if_stmt_992_branch_req_0 : boolean;
  signal addr_of_1156_final_reg_req_1 : boolean;
  signal if_stmt_992_branch_ack_1 : boolean;
  signal if_stmt_1239_branch_req_0 : boolean;
  signal if_stmt_992_branch_ack_0 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal type_cast_1002_inst_req_0 : boolean;
  signal type_cast_1002_inst_ack_0 : boolean;
  signal type_cast_1002_inst_req_1 : boolean;
  signal type_cast_1002_inst_ack_1 : boolean;
  signal type_cast_1258_inst_ack_1 : boolean;
  signal phi_stmt_902_req_1 : boolean;
  signal type_cast_1007_inst_req_0 : boolean;
  signal type_cast_1007_inst_ack_0 : boolean;
  signal type_cast_1007_inst_req_1 : boolean;
  signal type_cast_1007_inst_ack_1 : boolean;
  signal type_cast_1256_inst_ack_0 : boolean;
  signal phi_stmt_917_ack_0 : boolean;
  signal phi_stmt_910_ack_0 : boolean;
  signal type_cast_1041_inst_req_0 : boolean;
  signal type_cast_1232_inst_ack_1 : boolean;
  signal type_cast_1041_inst_ack_0 : boolean;
  signal phi_stmt_902_ack_0 : boolean;
  signal type_cast_1041_inst_req_1 : boolean;
  signal type_cast_1232_inst_req_1 : boolean;
  signal type_cast_1041_inst_ack_1 : boolean;
  signal type_cast_1258_inst_req_1 : boolean;
  signal phi_stmt_1246_req_1 : boolean;
  signal phi_stmt_917_req_0 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal phi_stmt_910_req_0 : boolean;
  signal type_cast_1149_inst_req_0 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal array_obj_ref_1047_index_offset_req_0 : boolean;
  signal array_obj_ref_1047_index_offset_ack_0 : boolean;
  signal array_obj_ref_1047_index_offset_req_1 : boolean;
  signal array_obj_ref_1047_index_offset_ack_1 : boolean;
  signal type_cast_1232_inst_ack_0 : boolean;
  signal type_cast_1232_inst_req_0 : boolean;
  signal addr_of_1048_final_reg_req_0 : boolean;
  signal addr_of_1048_final_reg_ack_0 : boolean;
  signal phi_stmt_917_req_1 : boolean;
  signal addr_of_1048_final_reg_req_1 : boolean;
  signal addr_of_1048_final_reg_ack_1 : boolean;
  signal phi_stmt_902_req_0 : boolean;
  signal type_cast_909_inst_ack_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal ptr_deref_1051_store_0_req_0 : boolean;
  signal ptr_deref_1159_store_0_ack_1 : boolean;
  signal ptr_deref_1051_store_0_ack_0 : boolean;
  signal ptr_deref_1051_store_0_req_1 : boolean;
  signal ptr_deref_1159_store_0_req_1 : boolean;
  signal ptr_deref_1051_store_0_ack_1 : boolean;
  signal type_cast_909_inst_req_1 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_1060_inst_req_0 : boolean;
  signal type_cast_1215_inst_ack_1 : boolean;
  signal type_cast_1060_inst_ack_0 : boolean;
  signal type_cast_1060_inst_req_1 : boolean;
  signal type_cast_1215_inst_req_1 : boolean;
  signal type_cast_1060_inst_ack_1 : boolean;
  signal addr_of_1156_final_reg_ack_0 : boolean;
  signal addr_of_1156_final_reg_req_0 : boolean;
  signal type_cast_1124_inst_req_0 : boolean;
  signal type_cast_1124_inst_ack_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal type_cast_1124_inst_req_1 : boolean;
  signal type_cast_1215_inst_ack_0 : boolean;
  signal type_cast_1124_inst_ack_1 : boolean;
  signal ptr_deref_1159_store_0_ack_0 : boolean;
  signal ptr_deref_1159_store_0_req_0 : boolean;
  signal type_cast_1258_inst_ack_0 : boolean;
  signal array_obj_ref_1130_index_offset_req_0 : boolean;
  signal array_obj_ref_1130_index_offset_ack_0 : boolean;
  signal array_obj_ref_1130_index_offset_req_1 : boolean;
  signal array_obj_ref_1130_index_offset_ack_1 : boolean;
  signal addr_of_1131_final_reg_req_0 : boolean;
  signal addr_of_1131_final_reg_ack_0 : boolean;
  signal addr_of_1131_final_reg_req_1 : boolean;
  signal addr_of_1131_final_reg_ack_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal ptr_deref_1135_load_0_req_0 : boolean;
  signal ptr_deref_1135_load_0_ack_0 : boolean;
  signal ptr_deref_1135_load_0_req_1 : boolean;
  signal ptr_deref_1135_load_0_ack_1 : boolean;
  signal phi_stmt_1246_ack_0 : boolean;
  signal phi_stmt_1253_ack_0 : boolean;
  signal phi_stmt_1259_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_A_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_A_CP_2408_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_A_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2408_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2408_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2408_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_A_CP_2408: Block -- control-path 
    signal zeropad3D_A_CP_2408_elements: BooleanArray(130 downto 0);
    -- 
  begin -- 
    zeropad3D_A_CP_2408_elements(0) <= zeropad3D_A_CP_2408_start;
    zeropad3D_A_CP_2408_symbol <= zeropad3D_A_CP_2408_elements(86);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_771/$entry
      -- CP-element group 0: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/$entry
      -- CP-element group 0: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_771/branch_block_stmt_771__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792__entry__
      -- 
    rr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(0), ack => RPIPE_Block0_starting_773_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	130 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	94 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	97 
    -- CP-element group 1: 	98 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_771/merge_stmt_1245__exit__
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Sample/rr
      -- 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(1), ack => type_cast_909_inst_req_0); -- 
    rr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(1), ack => type_cast_916_inst_req_0); -- 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(1), ack => type_cast_909_inst_req_1); -- 
    cr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(1), ack => type_cast_916_inst_req_1); -- 
    cr_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(1), ack => type_cast_923_inst_req_1); -- 
    rr_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(1), ack => type_cast_923_inst_req_0); -- 
    zeropad3D_A_CP_2408_elements(1) <= zeropad3D_A_CP_2408_elements(130);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_update_start_
      -- CP-element group 2: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Update/cr
      -- 
    ra_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_773_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(2)); -- 
    cr_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(2), ack => RPIPE_Block0_starting_773_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_773_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Sample/$entry
      -- 
    ca_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_773_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(3)); -- 
    rr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(3), ack => RPIPE_Block0_starting_776_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_update_start_
      -- CP-element group 4: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Update/cr
      -- 
    ra_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_776_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(4)); -- 
    cr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(4), ack => RPIPE_Block0_starting_776_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_776_Update/$exit
      -- 
    ca_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_776_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(5)); -- 
    rr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(5), ack => RPIPE_Block0_starting_779_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_update_start_
      -- CP-element group 6: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_sample_completed_
      -- 
    ra_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_779_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(6)); -- 
    cr_2507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(6), ack => RPIPE_Block0_starting_779_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_779_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Sample/rr
      -- 
    ca_2508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_779_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(7)); -- 
    rr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(7), ack => RPIPE_Block0_starting_782_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_update_start_
      -- CP-element group 8: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Update/cr
      -- 
    ra_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_782_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(8)); -- 
    cr_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(8), ack => RPIPE_Block0_starting_782_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_782_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Sample/rr
      -- 
    ca_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_782_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(9)); -- 
    rr_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(9), ack => RPIPE_Block0_starting_785_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_update_start_
      -- CP-element group 10: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Update/cr
      -- 
    ra_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_785_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(10)); -- 
    cr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(10), ack => RPIPE_Block0_starting_785_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_785_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Sample/rr
      -- 
    ca_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_785_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(11)); -- 
    rr_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(11), ack => RPIPE_Block0_starting_788_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_update_start_
      -- CP-element group 12: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Update/cr
      -- 
    ra_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_788_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(12)); -- 
    cr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(12), ack => RPIPE_Block0_starting_788_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_788_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Sample/rr
      -- 
    ca_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_788_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(13)); -- 
    rr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(13), ack => RPIPE_Block0_starting_791_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_update_start_
      -- CP-element group 14: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Update/cr
      -- 
    ra_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_791_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(14)); -- 
    cr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(14), ack => RPIPE_Block0_starting_791_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15:  members (49) 
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792__exit__
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/$exit
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899__entry__
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_774_to_assign_stmt_792/RPIPE_Block0_starting_791_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_update_start_
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Update/cr
      -- 
    ca_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_791_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(15)); -- 
    rr_2575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_796_inst_req_0); -- 
    cr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_796_inst_req_1); -- 
    rr_2589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_800_inst_req_0); -- 
    cr_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_800_inst_req_1); -- 
    rr_2603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_804_inst_req_0); -- 
    cr_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_804_inst_req_1); -- 
    rr_2617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_808_inst_req_0); -- 
    cr_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_808_inst_req_1); -- 
    rr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_817_inst_req_0); -- 
    cr_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_817_inst_req_1); -- 
    rr_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_821_inst_req_0); -- 
    cr_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_821_inst_req_1); -- 
    rr_2659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_857_inst_req_0); -- 
    cr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(15), ack => type_cast_857_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Sample/ra
      -- 
    ra_2576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_796_Update/ca
      -- 
    ca_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Sample/ra
      -- 
    ra_2590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	30 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_800_Update/ca
      -- 
    ca_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Sample/ra
      -- 
    ra_2604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	30 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_804_Update/ca
      -- 
    ca_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Sample/ra
      -- 
    ra_2618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_808_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	30 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_808_Update/ca
      -- 
    ca_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_808_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Sample/ra
      -- 
    ra_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_817_Update/ca
      -- 
    ca_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Sample/ra
      -- 
    ra_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_821_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_821_Update/ca
      -- 
    ca_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_821_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Sample/ra
      -- 
    ra_2660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/type_cast_857_Update/ca
      -- 
    ca_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: 	19 
    -- CP-element group 30: 	21 
    -- CP-element group 30: 	23 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	27 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	87 
    -- CP-element group 30: 	88 
    -- CP-element group 30: 	89 
    -- CP-element group 30:  members (10) 
      -- CP-element group 30: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899__exit__
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_771/assign_stmt_797_to_assign_stmt_899/$exit
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/$entry
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_917/$entry
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/$entry
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_910/$entry
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/$entry
      -- CP-element group 30: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_902/$entry
      -- 
    zeropad3D_A_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(17) & zeropad3D_A_CP_2408_elements(19) & zeropad3D_A_CP_2408_elements(21) & zeropad3D_A_CP_2408_elements(23) & zeropad3D_A_CP_2408_elements(25) & zeropad3D_A_CP_2408_elements(27) & zeropad3D_A_CP_2408_elements(29);
      gj_zeropad3D_A_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	105 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Sample/ra
      -- 
    ra_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(31)); -- 
    -- CP-element group 32:  branch  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	105 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (13) 
      -- CP-element group 32: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954__exit__
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955__entry__
      -- CP-element group 32: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/$exit
      -- CP-element group 32: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955_dead_link/$entry
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955_eval_test/$entry
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955_eval_test/$exit
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955_eval_test/branch_req
      -- CP-element group 32: 	 branch_block_stmt_771/R_orx_xcond_956_place
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955_if_link/$entry
      -- CP-element group 32: 	 branch_block_stmt_771/if_stmt_955_else_link/$entry
      -- 
    ca_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(32)); -- 
    branch_req_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(32), ack => if_stmt_955_branch_req_0); -- 
    -- CP-element group 33:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (18) 
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991__entry__
      -- CP-element group 33: 	 branch_block_stmt_771/merge_stmt_961__exit__
      -- CP-element group 33: 	 branch_block_stmt_771/merge_stmt_961_PhiAck/dummy
      -- CP-element group 33: 	 branch_block_stmt_771/merge_stmt_961_PhiReqMerge
      -- CP-element group 33: 	 branch_block_stmt_771/if_stmt_955_if_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_771/if_stmt_955_if_link/if_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_771/whilex_xbody_lorx_xlhsx_xfalse54
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/$entry
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_update_start_
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_771/merge_stmt_961_PhiAck/$exit
      -- CP-element group 33: 	 branch_block_stmt_771/merge_stmt_961_PhiAck/$entry
      -- CP-element group 33: 	 branch_block_stmt_771/whilex_xbody_lorx_xlhsx_xfalse54_PhiReq/$exit
      -- CP-element group 33: 	 branch_block_stmt_771/whilex_xbody_lorx_xlhsx_xfalse54_PhiReq/$entry
      -- 
    if_choice_transition_2695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_955_branch_ack_1, ack => zeropad3D_A_CP_2408_elements(33)); -- 
    rr_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(33), ack => type_cast_965_inst_req_0); -- 
    cr_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(33), ack => type_cast_965_inst_req_1); -- 
    -- CP-element group 34:  transition  place  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	106 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_771/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_771/if_stmt_955_else_link/$exit
      -- CP-element group 34: 	 branch_block_stmt_771/if_stmt_955_else_link/else_choice_transition
      -- CP-element group 34: 	 branch_block_stmt_771/whilex_xbody_ifx_xthen
      -- CP-element group 34: 	 branch_block_stmt_771/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_2699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_955_branch_ack_0, ack => zeropad3D_A_CP_2408_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Sample/ra
      -- 
    ra_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_965_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (13) 
      -- CP-element group 36: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991__exit__
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992__entry__
      -- CP-element group 36: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/$exit
      -- CP-element group 36: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_771/assign_stmt_966_to_assign_stmt_991/type_cast_965_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_771/R_orx_xcond186_993_place
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_771/if_stmt_992_else_link/$entry
      -- 
    ca_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_965_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(36)); -- 
    branch_req_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(36), ack => if_stmt_992_branch_req_0); -- 
    -- CP-element group 37:  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	71 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	68 
    -- CP-element group 37: 	64 
    -- CP-element group 37: 	53 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	56 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	60 
    -- CP-element group 37: 	62 
    -- CP-element group 37:  members (46) 
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161__entry__
      -- CP-element group 37: 	 branch_block_stmt_771/merge_stmt_1056_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/merge_stmt_1056_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_771/merge_stmt_1056_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_771/merge_stmt_1056__exit__
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_update_start_
      -- CP-element group 37: 	 branch_block_stmt_771/lorx_xlhsx_xfalse54_ifx_xelse_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_771/lorx_xlhsx_xfalse54_ifx_xelse_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_update_start
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_771/merge_stmt_1056_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_update_start_
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Update/req
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_complete/req
      -- CP-element group 37: 	 branch_block_stmt_771/if_stmt_992_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_771/if_stmt_992_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_771/lorx_xlhsx_xfalse54_ifx_xelse
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_update_start_
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_update_start_
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_update_start_
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_update_start
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Update/req
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_complete/req
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_update_start_
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_update_start_
      -- 
    if_choice_transition_2731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_992_branch_ack_1, ack => zeropad3D_A_CP_2408_elements(37)); -- 
    cr_3018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => type_cast_1149_inst_req_1); -- 
    req_3049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => array_obj_ref_1155_index_offset_req_1); -- 
    req_3064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => addr_of_1156_final_reg_req_1); -- 
    cr_3114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => ptr_deref_1159_store_0_req_1); -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => type_cast_1060_inst_req_0); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => type_cast_1060_inst_req_1); -- 
    cr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => type_cast_1124_inst_req_1); -- 
    req_2939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => array_obj_ref_1130_index_offset_req_1); -- 
    req_2954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => addr_of_1131_final_reg_req_1); -- 
    cr_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(37), ack => ptr_deref_1135_load_0_req_1); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	106 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_771/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_771/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$exit
      -- CP-element group 38: 	 branch_block_stmt_771/if_stmt_992_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_771/if_stmt_992_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_771/lorx_xlhsx_xfalse54_ifx_xthen
      -- 
    else_choice_transition_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_992_branch_ack_0, ack => zeropad3D_A_CP_2408_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	106 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Sample/ra
      -- 
    ra_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1002_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	106 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Update/ca
      -- 
    ca_2754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1002_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	106 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Sample/ra
      -- 
    ra_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1007_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	106 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Update/ca
      -- 
    ca_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1007_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Sample/rr
      -- 
    rr_2776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(43), ack => type_cast_1041_inst_req_0); -- 
    zeropad3D_A_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(40) & zeropad3D_A_CP_2408_elements(42);
      gj_zeropad3D_A_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Sample/ra
      -- 
    ra_2777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1041_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	106 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Sample/req
      -- 
    ca_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1041_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(45)); -- 
    req_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(45), ack => array_obj_ref_1047_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	52 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Sample/ack
      -- 
    ack_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1047_index_offset_ack_0, ack => zeropad3D_A_CP_2408_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	106 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_request/req
      -- 
    ack_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1047_index_offset_ack_1, ack => zeropad3D_A_CP_2408_elements(47)); -- 
    req_2822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(47), ack => addr_of_1048_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_request/ack
      -- 
    ack_2823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1048_final_reg_ack_0, ack => zeropad3D_A_CP_2408_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	106 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (28) 
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/ptr_deref_1051_Split/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/ptr_deref_1051_Split/$exit
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/ptr_deref_1051_Split/split_req
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/ptr_deref_1051_Split/split_ack
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/word_access_start/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/word_access_start/word_0/$entry
      -- CP-element group 49: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/word_access_start/word_0/rr
      -- 
    ack_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1048_final_reg_ack_1, ack => zeropad3D_A_CP_2408_elements(49)); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(49), ack => ptr_deref_1051_store_0_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Sample/word_access_start/word_0/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_store_0_ack_0, ack => zeropad3D_A_CP_2408_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	106 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/word_access_complete/word_0/ca
      -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_store_0_ack_1, ack => zeropad3D_A_CP_2408_elements(51)); -- 
    -- CP-element group 52:  join  transition  place  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	46 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	107 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_771/ifx_xthen_ifx_xend
      -- CP-element group 52: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054__exit__
      -- CP-element group 52: 	 branch_block_stmt_771/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_771/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/$exit
      -- 
    zeropad3D_A_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(46) & zeropad3D_A_CP_2408_elements(51);
      gj_zeropad3D_A_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	37 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Sample/ra
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1060_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	63 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1060_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_sample_start_
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1060_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(54)); -- 
    rr_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(54), ack => type_cast_1149_inst_req_0); -- 
    rr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(54), ack => type_cast_1124_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Sample/ra
      -- 
    ra_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1124_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	37 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (16) 
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1124_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Sample/req
      -- 
    ca_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1124_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(56)); -- 
    req_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(56), ack => array_obj_ref_1130_index_offset_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	72 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Sample/ack
      -- 
    ack_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1130_index_offset_ack_0, ack => zeropad3D_A_CP_2408_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1130_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_request/req
      -- 
    ack_2940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1130_index_offset_ack_1, ack => zeropad3D_A_CP_2408_elements(58)); -- 
    req_2949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(58), ack => addr_of_1131_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_request/ack
      -- 
    ack_2950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1131_final_reg_ack_0, ack => zeropad3D_A_CP_2408_elements(59)); -- 
    -- CP-element group 60:  join  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	37 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1131_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_word_addrgen/root_register_ack
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/word_access_start/$entry
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/word_access_start/word_0/$entry
      -- CP-element group 60: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/word_access_start/word_0/rr
      -- 
    ack_2955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1131_final_reg_ack_1, ack => zeropad3D_A_CP_2408_elements(60)); -- 
    rr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(60), ack => ptr_deref_1135_load_0_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/word_access_start/$exit
      -- CP-element group 61: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/word_access_start/word_0/$exit
      -- CP-element group 61: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Sample/word_access_start/word_0/ra
      -- 
    ra_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_load_0_ack_0, ack => zeropad3D_A_CP_2408_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	69 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/word_access_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/word_access_complete/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/word_access_complete/word_0/ca
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/ptr_deref_1135_Merge/$entry
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/ptr_deref_1135_Merge/$exit
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/ptr_deref_1135_Merge/merge_req
      -- CP-element group 62: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1135_Update/ptr_deref_1135_Merge/merge_ack
      -- 
    ca_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_load_0_ack_1, ack => zeropad3D_A_CP_2408_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	54 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_sample_completed_
      -- 
    ra_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	37 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (16) 
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_resized_1
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_scaled_1
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_computed_1
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_resize_1/$entry
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_resize_1/$exit
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_resize_1/index_resize_req
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_resize_1/index_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_scale_1/scale_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_scale_1/scale_rename_req
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_scale_1/$exit
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_index_scale_1/$entry
      -- CP-element group 64: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/type_cast_1149_update_completed_
      -- 
    ca_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(64)); -- 
    req_3044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(64), ack => array_obj_ref_1155_index_offset_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	72 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_sample_complete
      -- 
    ack_3045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1155_index_offset_ack_0, ack => zeropad3D_A_CP_2408_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (11) 
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_base_plus_offset/sum_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_offset_calculated
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_base_plus_offset/sum_rename_req
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_root_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_final_index_sum_regn_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_base_plus_offset/$entry
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/array_obj_ref_1155_base_plus_offset/$exit
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_request/req
      -- CP-element group 66: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_request/$entry
      -- 
    ack_3050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1155_index_offset_ack_1, ack => zeropad3D_A_CP_2408_elements(66)); -- 
    req_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(66), ack => addr_of_1156_final_reg_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_request/ack
      -- CP-element group 67: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_request/$exit
      -- 
    ack_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1156_final_reg_ack_0, ack => zeropad3D_A_CP_2408_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	37 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (19) 
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_address_resized
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_word_addrgen/$entry
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_addr_resize/$exit
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_word_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_addr_resize/base_resize_req
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_complete/ack
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_addr_resize/$entry
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_addr_resize/base_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/addr_of_1156_complete/$exit
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_word_addrgen/root_register_ack
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_word_addrgen/root_register_req
      -- CP-element group 68: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_word_addrgen/$exit
      -- 
    ack_3065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1156_final_reg_ack_1, ack => zeropad3D_A_CP_2408_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: 	62 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (9) 
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/ptr_deref_1159_Split/$exit
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/ptr_deref_1159_Split/$entry
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/word_access_start/word_0/rr
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/word_access_start/word_0/$entry
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/word_access_start/$entry
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/ptr_deref_1159_Split/split_ack
      -- CP-element group 69: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/ptr_deref_1159_Split/split_req
      -- 
    rr_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(69), ack => ptr_deref_1159_store_0_req_0); -- 
    zeropad3D_A_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(68) & zeropad3D_A_CP_2408_elements(62);
      gj_zeropad3D_A_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/word_access_start/word_0/ra
      -- CP-element group 70: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/word_access_start/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Sample/word_access_start/$exit
      -- 
    ra_3104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1159_store_0_ack_0, ack => zeropad3D_A_CP_2408_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	37 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/word_access_complete/word_0/ca
      -- CP-element group 71: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/word_access_complete/word_0/$exit
      -- CP-element group 71: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/word_access_complete/$exit
      -- CP-element group 71: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/ptr_deref_1159_Update/$exit
      -- 
    ca_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1159_store_0_ack_1, ack => zeropad3D_A_CP_2408_elements(71)); -- 
    -- CP-element group 72:  join  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: 	65 
    -- CP-element group 72: 	57 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	107 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_771/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_771/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_771/ifx_xelse_ifx_xend
      -- CP-element group 72: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161__exit__
      -- CP-element group 72: 	 branch_block_stmt_771/assign_stmt_1061_to_assign_stmt_1161/$exit
      -- 
    zeropad3D_A_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(71) & zeropad3D_A_CP_2408_elements(65) & zeropad3D_A_CP_2408_elements(57);
      gj_zeropad3D_A_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	107 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_sample_completed_
      -- 
    ra_3127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	107 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182__entry__
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181__exit__
      -- CP-element group 74: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_771/if_stmt_1182_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/$exit
      -- CP-element group 74: 	 branch_block_stmt_771/R_cmp139_1183_place
      -- 
    ca_3132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(74)); -- 
    branch_req_3140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(74), ack => if_stmt_1182_branch_req_0); -- 
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	116 
    -- CP-element group 75: 	117 
    -- CP-element group 75: 	119 
    -- CP-element group 75: 	120 
    -- CP-element group 75: 	122 
    -- CP-element group 75: 	123 
    -- CP-element group 75:  members (40) 
      -- CP-element group 75: 	 branch_block_stmt_771/merge_stmt_1188__exit__
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xend_ifx_xthen141_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/assign_stmt_1194__exit__
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180
      -- CP-element group 75: 	 branch_block_stmt_771/if_stmt_1182_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_771/merge_stmt_1188_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_771/merge_stmt_1188_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_771/merge_stmt_1188_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xend_ifx_xthen141_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_771/merge_stmt_1188_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_771/if_stmt_1182_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/assign_stmt_1194__entry__
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/assign_stmt_1194/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/assign_stmt_1194/$exit
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xend_ifx_xthen141
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/$entry
      -- CP-element group 75: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Sample/$entry
      -- 
    if_choice_transition_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1182_branch_ack_1, ack => zeropad3D_A_CP_2408_elements(75)); -- 
    cr_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(75), ack => type_cast_1256_inst_req_1); -- 
    rr_3487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(75), ack => type_cast_1249_inst_req_0); -- 
    rr_3533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(75), ack => type_cast_1262_inst_req_0); -- 
    cr_3538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(75), ack => type_cast_1262_inst_req_1); -- 
    cr_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(75), ack => type_cast_1249_inst_req_1); -- 
    rr_3510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(75), ack => type_cast_1256_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76: 	80 
    -- CP-element group 76: 	82 
    -- CP-element group 76:  members (24) 
      -- CP-element group 76: 	 branch_block_stmt_771/ifx_xend_ifx_xelse146
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238__entry__
      -- CP-element group 76: 	 branch_block_stmt_771/merge_stmt_1196__exit__
      -- CP-element group 76: 	 branch_block_stmt_771/if_stmt_1182_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_771/ifx_xend_ifx_xelse146_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_771/merge_stmt_1196_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_771/ifx_xend_ifx_xelse146_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_771/if_stmt_1182_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_771/merge_stmt_1196_PhiAck/$entry
      -- CP-element group 76: 	 branch_block_stmt_771/merge_stmt_1196_PhiAck/$exit
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_771/merge_stmt_1196_PhiAck/dummy
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_update_start_
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_update_start_
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_update_start_
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/$entry
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Update/$entry
      -- 
    else_choice_transition_3149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1182_branch_ack_0, ack => zeropad3D_A_CP_2408_elements(76)); -- 
    rr_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(76), ack => type_cast_1206_inst_req_0); -- 
    cr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(76), ack => type_cast_1206_inst_req_1); -- 
    cr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(76), ack => type_cast_1232_inst_req_1); -- 
    cr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(76), ack => type_cast_1215_inst_req_1); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_sample_completed_
      -- 
    ra_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1206_update_completed_
      -- 
    ca_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(78)); -- 
    rr_3179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(78), ack => type_cast_1215_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Sample/ra
      -- 
    ra_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	76 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1215_Update/$exit
      -- 
    ca_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(80)); -- 
    rr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(80), ack => type_cast_1232_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_sample_completed_
      -- 
    ra_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1232_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(81)); -- 
    -- CP-element group 82:  branch  transition  place  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	76 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (13) 
      -- CP-element group 82: 	 branch_block_stmt_771/R_cmp172_1240_place
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239__entry__
      -- CP-element group 82: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238__exit__
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239_if_link/$entry
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239_else_link/$entry
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239_eval_test/branch_req
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239_eval_test/$exit
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239_eval_test/$entry
      -- CP-element group 82: 	 branch_block_stmt_771/if_stmt_1239_dead_link/$entry
      -- CP-element group 82: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/type_cast_1232_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_771/assign_stmt_1202_to_assign_stmt_1238/$exit
      -- 
    ca_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1232_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(82)); -- 
    branch_req_3207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(82), ack => if_stmt_1239_branch_req_0); -- 
    -- CP-element group 83:  transition  place  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (15) 
      -- CP-element group 83: 	 branch_block_stmt_771/merge_stmt_1267__exit__
      -- CP-element group 83: 	 branch_block_stmt_771/assign_stmt_1272__entry__
      -- CP-element group 83: 	 branch_block_stmt_771/ifx_xelse146_whilex_xend
      -- CP-element group 83: 	 branch_block_stmt_771/if_stmt_1239_if_link/if_choice_transition
      -- CP-element group 83: 	 branch_block_stmt_771/if_stmt_1239_if_link/$exit
      -- CP-element group 83: 	 branch_block_stmt_771/assign_stmt_1272/$entry
      -- CP-element group 83: 	 branch_block_stmt_771/merge_stmt_1267_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Sample/req
      -- CP-element group 83: 	 branch_block_stmt_771/ifx_xelse146_whilex_xend_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_771/ifx_xelse146_whilex_xend_PhiReq/$exit
      -- CP-element group 83: 	 branch_block_stmt_771/merge_stmt_1267_PhiAck/$entry
      -- CP-element group 83: 	 branch_block_stmt_771/merge_stmt_1267_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_771/merge_stmt_1267_PhiAck/dummy
      -- 
    if_choice_transition_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1239_branch_ack_1, ack => zeropad3D_A_CP_2408_elements(83)); -- 
    req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(83), ack => WPIPE_Block0_complete_1269_inst_req_0); -- 
    -- CP-element group 84:  fork  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	108 
    -- CP-element group 84: 	109 
    -- CP-element group 84: 	110 
    -- CP-element group 84: 	112 
    -- CP-element group 84: 	113 
    -- CP-element group 84:  members (22) 
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180
      -- CP-element group 84: 	 branch_block_stmt_771/if_stmt_1239_else_link/$exit
      -- CP-element group 84: 	 branch_block_stmt_771/if_stmt_1239_else_link/else_choice_transition
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Update/cr
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1246/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Update/cr
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/$entry
      -- 
    else_choice_transition_3216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1239_branch_ack_0, ack => zeropad3D_A_CP_2408_elements(84)); -- 
    rr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(84), ack => type_cast_1264_inst_req_0); -- 
    cr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(84), ack => type_cast_1264_inst_req_1); -- 
    rr_3438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(84), ack => type_cast_1258_inst_req_0); -- 
    cr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(84), ack => type_cast_1258_inst_req_1); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_update_start_
      -- CP-element group 85: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Sample/ack
      -- CP-element group 85: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Update/req
      -- 
    ack_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1269_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(85)); -- 
    req_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(85), ack => WPIPE_Block0_complete_1269_inst_req_1); -- 
    -- CP-element group 86:  transition  place  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_771/return__
      -- CP-element group 86: 	 branch_block_stmt_771/assign_stmt_1272__exit__
      -- CP-element group 86: 	 $exit
      -- CP-element group 86: 	 branch_block_stmt_771/merge_stmt_1274__exit__
      -- CP-element group 86: 	 branch_block_stmt_771/$exit
      -- CP-element group 86: 	 branch_block_stmt_771/branch_block_stmt_771__exit__
      -- CP-element group 86: 	 branch_block_stmt_771/assign_stmt_1272/$exit
      -- CP-element group 86: 	 branch_block_stmt_771/merge_stmt_1274_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_771/assign_stmt_1272/WPIPE_Block0_complete_1269_Update/ack
      -- CP-element group 86: 	 branch_block_stmt_771/return___PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_771/return___PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_771/merge_stmt_1274_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_771/merge_stmt_1274_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_771/merge_stmt_1274_PhiAck/dummy
      -- 
    ack_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1269_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(86)); -- 
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	30 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_req
      -- CP-element group 87: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_907_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_902/$exit
      -- 
    phi_stmt_902_req_3246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_902_req_3246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(87), ack => phi_stmt_902_req_0); -- 
    -- Element group zeropad3D_A_CP_2408_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2408_elements(30), ack => zeropad3D_A_CP_2408_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  transition  output  delay-element  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	30 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_req
      -- CP-element group 88: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_914_konst_delay_trans
      -- CP-element group 88: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_910/$exit
      -- 
    phi_stmt_910_req_3254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_910_req_3254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(88), ack => phi_stmt_910_req_0); -- 
    -- Element group zeropad3D_A_CP_2408_elements(88) is a control-delay.
    cp_element_88_delay: control_delay_element  generic map(name => " 88_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2408_elements(30), ack => zeropad3D_A_CP_2408_elements(88), clk => clk, reset =>reset);
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	30 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_req
      -- CP-element group 89: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_921_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/phi_stmt_917/$exit
      -- 
    phi_stmt_917_req_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_917_req_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(89), ack => phi_stmt_917_req_0); -- 
    -- Element group zeropad3D_A_CP_2408_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2408_elements(30), ack => zeropad3D_A_CP_2408_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  join  transition  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	101 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_771/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(87) & zeropad3D_A_CP_2408_elements(88) & zeropad3D_A_CP_2408_elements(89);
      gj_zeropad3D_A_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Sample/ra
      -- 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_909_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Update/ca
      -- CP-element group 92: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/Update/$exit
      -- 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_909_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	100 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/type_cast_909/$exit
      -- CP-element group 93: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/phi_stmt_902_req
      -- CP-element group 93: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_902/$exit
      -- 
    phi_stmt_902_req_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_902_req_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(93), ack => phi_stmt_902_req_1); -- 
    zeropad3D_A_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(91) & zeropad3D_A_CP_2408_elements(92);
      gj_zeropad3D_A_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Sample/ra
      -- 
    ra_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/Update/ca
      -- 
    ca_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_req
      -- CP-element group 96: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/$exit
      -- CP-element group 96: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/$exit
      -- CP-element group 96: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_910/phi_stmt_910_sources/type_cast_916/SplitProtocol/$exit
      -- 
    phi_stmt_910_req_3311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_910_req_3311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(96), ack => phi_stmt_910_req_1); -- 
    zeropad3D_A_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(94) & zeropad3D_A_CP_2408_elements(95);
      gj_zeropad3D_A_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	1 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Sample/ra
      -- 
    ra_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Update/ca
      -- CP-element group 98: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/Update/$exit
      -- 
    ca_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/$exit
      -- CP-element group 99: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/$exit
      -- CP-element group 99: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_sources/type_cast_923/SplitProtocol/$exit
      -- CP-element group 99: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_917/phi_stmt_917_req
      -- 
    phi_stmt_917_req_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_917_req_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(99), ack => phi_stmt_917_req_1); -- 
    zeropad3D_A_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(97) & zeropad3D_A_CP_2408_elements(98);
      gj_zeropad3D_A_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	93 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_771/ifx_xend180_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(93) & zeropad3D_A_CP_2408_elements(96) & zeropad3D_A_CP_2408_elements(99);
      gj_zeropad3D_A_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  merge  fork  transition  place  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	90 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_771/merge_stmt_901_PhiReqMerge
      -- CP-element group 101: 	 branch_block_stmt_771/merge_stmt_901_PhiAck/$entry
      -- 
    zeropad3D_A_CP_2408_elements(101) <= OrReduce(zeropad3D_A_CP_2408_elements(90) & zeropad3D_A_CP_2408_elements(100));
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	105 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_771/merge_stmt_901_PhiAck/phi_stmt_902_ack
      -- 
    phi_stmt_902_ack_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_902_ack_0, ack => zeropad3D_A_CP_2408_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_771/merge_stmt_901_PhiAck/phi_stmt_910_ack
      -- 
    phi_stmt_910_ack_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_910_ack_0, ack => zeropad3D_A_CP_2408_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	101 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_771/merge_stmt_901_PhiAck/phi_stmt_917_ack
      -- 
    phi_stmt_917_ack_3341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_917_ack_0, ack => zeropad3D_A_CP_2408_elements(104)); -- 
    -- CP-element group 105:  join  fork  transition  place  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	102 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	31 
    -- CP-element group 105: 	32 
    -- CP-element group 105:  members (10) 
      -- CP-element group 105: 	 branch_block_stmt_771/merge_stmt_901__exit__
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954__entry__
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/$entry
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_update_start_
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_771/assign_stmt_929_to_assign_stmt_954/type_cast_928_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_771/merge_stmt_901_PhiAck/$exit
      -- 
    rr_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(105), ack => type_cast_928_inst_req_0); -- 
    cr_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(105), ack => type_cast_928_inst_req_1); -- 
    zeropad3D_A_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(102) & zeropad3D_A_CP_2408_elements(103) & zeropad3D_A_CP_2408_elements(104);
      gj_zeropad3D_A_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  merge  fork  transition  place  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	34 
    -- CP-element group 106: 	38 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	39 
    -- CP-element group 106: 	40 
    -- CP-element group 106: 	41 
    -- CP-element group 106: 	42 
    -- CP-element group 106: 	45 
    -- CP-element group 106: 	47 
    -- CP-element group 106: 	49 
    -- CP-element group 106: 	51 
    -- CP-element group 106:  members (33) 
      -- CP-element group 106: 	 branch_block_stmt_771/merge_stmt_998__exit__
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054__entry__
      -- CP-element group 106: 	 branch_block_stmt_771/merge_stmt_998_PhiReqMerge
      -- CP-element group 106: 	 branch_block_stmt_771/merge_stmt_998_PhiAck/dummy
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_update_start_
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1002_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_update_start_
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1007_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_update_start_
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/type_cast_1041_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_update_start_
      -- CP-element group 106: 	 branch_block_stmt_771/merge_stmt_998_PhiAck/$exit
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_update_start
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/array_obj_ref_1047_final_index_sum_regn_Update/req
      -- CP-element group 106: 	 branch_block_stmt_771/merge_stmt_998_PhiAck/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_complete/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/addr_of_1048_complete/req
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_update_start_
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/word_access_complete/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/word_access_complete/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_771/assign_stmt_1003_to_assign_stmt_1054/ptr_deref_1051_Update/word_access_complete/word_0/cr
      -- 
    rr_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => type_cast_1002_inst_req_0); -- 
    cr_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => type_cast_1002_inst_req_1); -- 
    rr_2762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => type_cast_1007_inst_req_0); -- 
    cr_2767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => type_cast_1007_inst_req_1); -- 
    cr_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => type_cast_1041_inst_req_1); -- 
    req_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => array_obj_ref_1047_index_offset_req_1); -- 
    req_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => addr_of_1048_final_reg_req_1); -- 
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(106), ack => ptr_deref_1051_store_0_req_1); -- 
    zeropad3D_A_CP_2408_elements(106) <= OrReduce(zeropad3D_A_CP_2408_elements(34) & zeropad3D_A_CP_2408_elements(38));
    -- CP-element group 107:  merge  fork  transition  place  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	72 
    -- CP-element group 107: 	52 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	73 
    -- CP-element group 107: 	74 
    -- CP-element group 107:  members (13) 
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_771/merge_stmt_1163__exit__
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181__entry__
      -- CP-element group 107: 	 branch_block_stmt_771/merge_stmt_1163_PhiAck/dummy
      -- CP-element group 107: 	 branch_block_stmt_771/merge_stmt_1163_PhiAck/$exit
      -- CP-element group 107: 	 branch_block_stmt_771/merge_stmt_1163_PhiAck/$entry
      -- CP-element group 107: 	 branch_block_stmt_771/merge_stmt_1163_PhiReqMerge
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_update_start_
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/type_cast_1167_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_771/assign_stmt_1168_to_assign_stmt_1181/$entry
      -- 
    cr_3131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(107), ack => type_cast_1167_inst_req_1); -- 
    rr_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(107), ack => type_cast_1167_inst_req_0); -- 
    zeropad3D_A_CP_2408_elements(107) <= OrReduce(zeropad3D_A_CP_2408_elements(72) & zeropad3D_A_CP_2408_elements(52));
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	84 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	115 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_req
      -- CP-element group 108: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1252_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1246/$exit
      -- 
    phi_stmt_1246_req_3422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1246_req_3422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(108), ack => phi_stmt_1246_req_1); -- 
    -- Element group zeropad3D_A_CP_2408_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2408_elements(84), ack => zeropad3D_A_CP_2408_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	84 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Sample/ra
      -- 
    ra_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	84 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Update/ca
      -- CP-element group 110: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/Update/$exit
      -- 
    ca_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	115 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/$exit
      -- CP-element group 111: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1258/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_req
      -- CP-element group 111: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1253/$exit
      -- 
    phi_stmt_1253_req_3445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1253_req_3445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(111), ack => phi_stmt_1253_req_1); -- 
    zeropad3D_A_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(109) & zeropad3D_A_CP_2408_elements(110);
      gj_zeropad3D_A_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	84 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Sample/ra
      -- 
    ra_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1264_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	84 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/Update/ca
      -- 
    ca_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1264_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/$exit
      -- CP-element group 114: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_req
      -- CP-element group 114: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1264/$exit
      -- CP-element group 114: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/$exit
      -- 
    phi_stmt_1259_req_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1259_req_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(114), ack => phi_stmt_1259_req_1); -- 
    zeropad3D_A_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(112) & zeropad3D_A_CP_2408_elements(113);
      gj_zeropad3D_A_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	108 
    -- CP-element group 115: 	111 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	126 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_771/ifx_xelse146_ifx_xend180_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(108) & zeropad3D_A_CP_2408_elements(111) & zeropad3D_A_CP_2408_elements(114);
      gj_zeropad3D_A_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	75 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Sample/$exit
      -- 
    ra_3488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	75 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/Update/$exit
      -- 
    ca_3493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	125 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/$exit
      -- CP-element group 118: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/$exit
      -- CP-element group 118: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_sources/type_cast_1249/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1246/phi_stmt_1246_req
      -- 
    phi_stmt_1246_req_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1246_req_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(118), ack => phi_stmt_1246_req_0); -- 
    zeropad3D_A_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(116) & zeropad3D_A_CP_2408_elements(117);
      gj_zeropad3D_A_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Sample/ra
      -- 
    ra_3511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	75 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/Update/$exit
      -- 
    ca_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	125 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/$exit
      -- CP-element group 121: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_req
      -- CP-element group 121: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1253/phi_stmt_1253_sources/type_cast_1256/$exit
      -- 
    phi_stmt_1253_req_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1253_req_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(121), ack => phi_stmt_1253_req_0); -- 
    zeropad3D_A_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(119) & zeropad3D_A_CP_2408_elements(120);
      gj_zeropad3D_A_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	75 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Sample/$exit
      -- 
    ra_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1262_inst_ack_0, ack => zeropad3D_A_CP_2408_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	75 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/Update/ca
      -- 
    ca_3539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1262_inst_ack_1, ack => zeropad3D_A_CP_2408_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/$exit
      -- CP-element group 124: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/$exit
      -- CP-element group 124: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_req
      -- CP-element group 124: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/$exit
      -- CP-element group 124: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1259/phi_stmt_1259_sources/type_cast_1262/SplitProtocol/$exit
      -- 
    phi_stmt_1259_req_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1259_req_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2408_elements(124), ack => phi_stmt_1259_req_0); -- 
    zeropad3D_A_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(122) & zeropad3D_A_CP_2408_elements(123);
      gj_zeropad3D_A_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	118 
    -- CP-element group 125: 	121 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_771/ifx_xthen141_ifx_xend180_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(118) & zeropad3D_A_CP_2408_elements(121) & zeropad3D_A_CP_2408_elements(124);
      gj_zeropad3D_A_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  merge  fork  transition  place  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	115 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126: 	129 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_771/merge_stmt_1245_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_771/merge_stmt_1245_PhiAck/$entry
      -- 
    zeropad3D_A_CP_2408_elements(126) <= OrReduce(zeropad3D_A_CP_2408_elements(115) & zeropad3D_A_CP_2408_elements(125));
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	130 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_771/merge_stmt_1245_PhiAck/phi_stmt_1246_ack
      -- 
    phi_stmt_1246_ack_3545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1246_ack_0, ack => zeropad3D_A_CP_2408_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_771/merge_stmt_1245_PhiAck/phi_stmt_1253_ack
      -- 
    phi_stmt_1253_ack_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1253_ack_0, ack => zeropad3D_A_CP_2408_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_771/merge_stmt_1245_PhiAck/phi_stmt_1259_ack
      -- 
    phi_stmt_1259_ack_3547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1259_ack_0, ack => zeropad3D_A_CP_2408_elements(129)); -- 
    -- CP-element group 130:  join  transition  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	127 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	1 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_771/merge_stmt_1245_PhiAck/$exit
      -- 
    zeropad3D_A_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2408_elements(127) & zeropad3D_A_CP_2408_elements(128) & zeropad3D_A_CP_2408_elements(129);
      gj_zeropad3D_A_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2408_elements(130), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1035_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1118_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1143_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_835_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_897_wire : std_logic_vector(31 downto 0);
    signal R_idxprom126_1129_resized : std_logic_vector(13 downto 0);
    signal R_idxprom126_1129_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom131_1154_resized : std_logic_vector(13 downto 0);
    signal R_idxprom131_1154_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1046_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1046_scaled : std_logic_vector(13 downto 0);
    signal add107_1091 : std_logic_vector(31 downto 0);
    signal add117_1106 : std_logic_vector(31 downto 0);
    signal add123_1111 : std_logic_vector(31 downto 0);
    signal add136_1174 : std_logic_vector(31 downto 0);
    signal add144_1194 : std_logic_vector(15 downto 0);
    signal add155_854 : std_logic_vector(31 downto 0);
    signal add171_869 : std_logic_vector(31 downto 0);
    signal add69_879 : std_logic_vector(31 downto 0);
    signal add80_1023 : std_logic_vector(31 downto 0);
    signal add86_1028 : std_logic_vector(31 downto 0);
    signal add98_1086 : std_logic_vector(31 downto 0);
    signal add_874 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1047_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1047_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1047_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1047_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1047_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1047_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1130_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1130_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1130_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1130_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1130_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1130_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_root_address : std_logic_vector(13 downto 0);
    signal arrayidx127_1132 : std_logic_vector(31 downto 0);
    signal arrayidx132_1157 : std_logic_vector(31 downto 0);
    signal arrayidx_1049 : std_logic_vector(31 downto 0);
    signal call1_777 : std_logic_vector(7 downto 0);
    signal call2_780 : std_logic_vector(7 downto 0);
    signal call3_783 : std_logic_vector(7 downto 0);
    signal call4_786 : std_logic_vector(7 downto 0);
    signal call5_789 : std_logic_vector(7 downto 0);
    signal call6_792 : std_logic_vector(7 downto 0);
    signal call_774 : std_logic_vector(7 downto 0);
    signal cmp139_1181 : std_logic_vector(0 downto 0);
    signal cmp156_1212 : std_logic_vector(0 downto 0);
    signal cmp172_1238 : std_logic_vector(0 downto 0);
    signal cmp52_949 : std_logic_vector(0 downto 0);
    signal cmp59_973 : std_logic_vector(0 downto 0);
    signal cmp59x_xnot_979 : std_logic_vector(0 downto 0);
    signal cmp70_986 : std_logic_vector(0 downto 0);
    signal cmp_936 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_942 : std_logic_vector(0 downto 0);
    signal conv100_899 : std_logic_vector(31 downto 0);
    signal conv135_1168 : std_logic_vector(31 downto 0);
    signal conv149_1207 : std_logic_vector(31 downto 0);
    signal conv164_1233 : std_logic_vector(31 downto 0);
    signal conv166_858 : std_logic_vector(31 downto 0);
    signal conv27_797 : std_logic_vector(31 downto 0);
    signal conv29_801 : std_logic_vector(31 downto 0);
    signal conv33_805 : std_logic_vector(31 downto 0);
    signal conv35_809 : std_logic_vector(31 downto 0);
    signal conv42_929 : std_logic_vector(31 downto 0);
    signal conv44_818 : std_logic_vector(31 downto 0);
    signal conv56_966 : std_logic_vector(31 downto 0);
    signal conv74_1003 : std_logic_vector(31 downto 0);
    signal conv76_822 : std_logic_vector(31 downto 0);
    signal conv78_1008 : std_logic_vector(31 downto 0);
    signal conv82_837 : std_logic_vector(31 downto 0);
    signal conv90_1061 : std_logic_vector(31 downto 0);
    signal div152_843 : std_logic_vector(31 downto 0);
    signal div167_864 : std_logic_vector(31 downto 0);
    signal idxprom126_1125 : std_logic_vector(63 downto 0);
    signal idxprom131_1150 : std_logic_vector(63 downto 0);
    signal idxprom_1042 : std_logic_vector(63 downto 0);
    signal inc161_1216 : std_logic_vector(15 downto 0);
    signal inc161x_xix_x2_1221 : std_logic_vector(15 downto 0);
    signal inc_1202 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1253 : std_logic_vector(15 downto 0);
    signal ix_x2_910 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1259 : std_logic_vector(15 downto 0);
    signal jx_x1_917 : std_logic_vector(15 downto 0);
    signal jx_x2_1228 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1246 : std_logic_vector(15 downto 0);
    signal kx_x1_902 : std_logic_vector(15 downto 0);
    signal mul106_1081 : std_logic_vector(31 downto 0);
    signal mul116_1096 : std_logic_vector(31 downto 0);
    signal mul122_1101 : std_logic_vector(31 downto 0);
    signal mul36_814 : std_logic_vector(31 downto 0);
    signal mul79_1013 : std_logic_vector(31 downto 0);
    signal mul85_1018 : std_logic_vector(31 downto 0);
    signal mul97_1071 : std_logic_vector(31 downto 0);
    signal mul_885 : std_logic_vector(31 downto 0);
    signal orx_xcond186_991 : std_logic_vector(0 downto 0);
    signal orx_xcond_954 : std_logic_vector(0 downto 0);
    signal ptr_deref_1051_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1051_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1051_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1051_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1051_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1051_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1135_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1135_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1135_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1135_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1135_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1159_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1159_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1159_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1159_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1159_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1159_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext185_828 : std_logic_vector(31 downto 0);
    signal sext_890 : std_logic_vector(31 downto 0);
    signal shl_849 : std_logic_vector(31 downto 0);
    signal shr125_1120 : std_logic_vector(31 downto 0);
    signal shr130_1145 : std_logic_vector(31 downto 0);
    signal shr_1037 : std_logic_vector(31 downto 0);
    signal sub105_1076 : std_logic_vector(31 downto 0);
    signal sub_1066 : std_logic_vector(31 downto 0);
    signal tmp128_1136 : std_logic_vector(63 downto 0);
    signal type_cast_1001_wire : std_logic_vector(31 downto 0);
    signal type_cast_1006_wire : std_logic_vector(31 downto 0);
    signal type_cast_1031_wire : std_logic_vector(31 downto 0);
    signal type_cast_1034_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1040_wire : std_logic_vector(63 downto 0);
    signal type_cast_1053_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1059_wire : std_logic_vector(31 downto 0);
    signal type_cast_1114_wire : std_logic_vector(31 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1123_wire : std_logic_vector(63 downto 0);
    signal type_cast_1139_wire : std_logic_vector(31 downto 0);
    signal type_cast_1142_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1148_wire : std_logic_vector(63 downto 0);
    signal type_cast_1166_wire : std_logic_vector(31 downto 0);
    signal type_cast_1172_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1177_wire : std_logic_vector(31 downto 0);
    signal type_cast_1179_wire : std_logic_vector(31 downto 0);
    signal type_cast_1192_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1200_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1205_wire : std_logic_vector(31 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1231_wire : std_logic_vector(31 downto 0);
    signal type_cast_1249_wire : std_logic_vector(15 downto 0);
    signal type_cast_1252_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1256_wire : std_logic_vector(15 downto 0);
    signal type_cast_1258_wire : std_logic_vector(15 downto 0);
    signal type_cast_1262_wire : std_logic_vector(15 downto 0);
    signal type_cast_1264_wire : std_logic_vector(15 downto 0);
    signal type_cast_1271_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_826_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_831_wire : std_logic_vector(31 downto 0);
    signal type_cast_834_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_841_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_847_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_862_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_883_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_893_wire : std_logic_vector(31 downto 0);
    signal type_cast_896_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_907_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_909_wire : std_logic_vector(15 downto 0);
    signal type_cast_914_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_916_wire : std_logic_vector(15 downto 0);
    signal type_cast_921_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_923_wire : std_logic_vector(15 downto 0);
    signal type_cast_927_wire : std_logic_vector(31 downto 0);
    signal type_cast_932_wire : std_logic_vector(31 downto 0);
    signal type_cast_934_wire : std_logic_vector(31 downto 0);
    signal type_cast_940_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_945_wire : std_logic_vector(31 downto 0);
    signal type_cast_947_wire : std_logic_vector(31 downto 0);
    signal type_cast_964_wire : std_logic_vector(31 downto 0);
    signal type_cast_969_wire : std_logic_vector(31 downto 0);
    signal type_cast_971_wire : std_logic_vector(31 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_982_wire : std_logic_vector(31 downto 0);
    signal type_cast_984_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1047_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1047_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1047_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1047_resized_base_address <= "00000000000000";
    array_obj_ref_1130_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1130_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1130_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1130_resized_base_address <= "00000000000000";
    array_obj_ref_1155_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1155_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1155_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1155_resized_base_address <= "00000000000000";
    ptr_deref_1051_word_offset_0 <= "00000000000000";
    ptr_deref_1135_word_offset_0 <= "00000000000000";
    ptr_deref_1159_word_offset_0 <= "00000000000000";
    type_cast_1034_wire_constant <= "00000000000000000000000000000010";
    type_cast_1053_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1117_wire_constant <= "00000000000000000000000000000010";
    type_cast_1142_wire_constant <= "00000000000000000000000000000010";
    type_cast_1172_wire_constant <= "00000000000000000000000000000100";
    type_cast_1192_wire_constant <= "0000000000000100";
    type_cast_1200_wire_constant <= "0000000000000001";
    type_cast_1225_wire_constant <= "0000000000000000";
    type_cast_1252_wire_constant <= "0000000000000000";
    type_cast_1271_wire_constant <= "00000001";
    type_cast_826_wire_constant <= "00000000000000000000000000010000";
    type_cast_834_wire_constant <= "00000000000000000000000000010000";
    type_cast_841_wire_constant <= "00000000000000000000000000000001";
    type_cast_847_wire_constant <= "00000000000000000000000000000001";
    type_cast_862_wire_constant <= "00000000000000000000000000000010";
    type_cast_883_wire_constant <= "00000000000000000000000000010000";
    type_cast_896_wire_constant <= "00000000000000000000000000010000";
    type_cast_907_wire_constant <= "0000000000000000";
    type_cast_914_wire_constant <= "0000000000000000";
    type_cast_921_wire_constant <= "0000000000000000";
    type_cast_940_wire_constant <= "1";
    type_cast_977_wire_constant <= "1";
    phi_stmt_1246: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1249_wire & type_cast_1252_wire_constant;
      req <= phi_stmt_1246_req_0 & phi_stmt_1246_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1246",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1246_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1246,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1246
    phi_stmt_1253: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1256_wire & type_cast_1258_wire;
      req <= phi_stmt_1253_req_0 & phi_stmt_1253_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1253",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1253_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1253,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1253
    phi_stmt_1259: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1262_wire & type_cast_1264_wire;
      req <= phi_stmt_1259_req_0 & phi_stmt_1259_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1259",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1259_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1259,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1259
    phi_stmt_902: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_907_wire_constant & type_cast_909_wire;
      req <= phi_stmt_902_req_0 & phi_stmt_902_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_902",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_902_ack_0,
          idata => idata,
          odata => kx_x1_902,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_902
    phi_stmt_910: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_914_wire_constant & type_cast_916_wire;
      req <= phi_stmt_910_req_0 & phi_stmt_910_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_910",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_910_ack_0,
          idata => idata,
          odata => ix_x2_910,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_910
    phi_stmt_917: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_921_wire_constant & type_cast_923_wire;
      req <= phi_stmt_917_req_0 & phi_stmt_917_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_917",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_917_ack_0,
          idata => idata,
          odata => jx_x1_917,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_917
    -- flow-through select operator MUX_1227_inst
    jx_x2_1228 <= type_cast_1225_wire_constant when (cmp156_1212(0) /=  '0') else inc_1202;
    addr_of_1048_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1048_final_reg_req_0;
      addr_of_1048_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1048_final_reg_req_1;
      addr_of_1048_final_reg_ack_1<= rack(0);
      addr_of_1048_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1048_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1047_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1131_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1131_final_reg_req_0;
      addr_of_1131_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1131_final_reg_req_1;
      addr_of_1131_final_reg_ack_1<= rack(0);
      addr_of_1131_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1131_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1130_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx127_1132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1156_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1156_final_reg_req_0;
      addr_of_1156_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1156_final_reg_req_1;
      addr_of_1156_final_reg_ack_1<= rack(0);
      addr_of_1156_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1156_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1155_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx132_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1002_inst_req_0;
      type_cast_1002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1002_inst_req_1;
      type_cast_1002_inst_ack_1<= rack(0);
      type_cast_1002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1002_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1001_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1007_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1007_inst_req_0;
      type_cast_1007_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1007_inst_req_1;
      type_cast_1007_inst_ack_1<= rack(0);
      type_cast_1007_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1007_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1006_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_1008,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1031_inst
    process(add86_1028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add86_1028(31 downto 0);
      type_cast_1031_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1036_inst
    process(ASHR_i32_i32_1035_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1035_wire(31 downto 0);
      shr_1037 <= tmp_var; -- 
    end process;
    type_cast_1041_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1041_inst_req_0;
      type_cast_1041_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1041_inst_req_1;
      type_cast_1041_inst_ack_1<= rack(0);
      type_cast_1041_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1041_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1040_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1042,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1060_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1060_inst_req_0;
      type_cast_1060_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1060_inst_req_1;
      type_cast_1060_inst_ack_1<= rack(0);
      type_cast_1060_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1060_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1059_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1061,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1114_inst
    process(add107_1091) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add107_1091(31 downto 0);
      type_cast_1114_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1119_inst
    process(ASHR_i32_i32_1118_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1118_wire(31 downto 0);
      shr125_1120 <= tmp_var; -- 
    end process;
    type_cast_1124_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1124_inst_req_0;
      type_cast_1124_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1124_inst_req_1;
      type_cast_1124_inst_ack_1<= rack(0);
      type_cast_1124_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1124_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1123_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom126_1125,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1139_inst
    process(add123_1111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add123_1111(31 downto 0);
      type_cast_1139_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1144_inst
    process(ASHR_i32_i32_1143_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1143_wire(31 downto 0);
      shr130_1145 <= tmp_var; -- 
    end process;
    type_cast_1149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1149_inst_req_0;
      type_cast_1149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1149_inst_req_1;
      type_cast_1149_inst_ack_1<= rack(0);
      type_cast_1149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1148_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom131_1150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1166_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1177_inst
    process(add136_1174) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add136_1174(31 downto 0);
      type_cast_1177_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1179_inst
    process(conv27_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv27_797(31 downto 0);
      type_cast_1179_wire <= tmp_var; -- 
    end process;
    type_cast_1206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1206_inst_req_0;
      type_cast_1206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1206_inst_req_1;
      type_cast_1206_inst_ack_1<= rack(0);
      type_cast_1206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1205_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_1207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1215_inst_req_0;
      type_cast_1215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1215_inst_req_1;
      type_cast_1215_inst_ack_1<= rack(0);
      type_cast_1215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp156_1212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc161_1216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1232_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1232_inst_req_0;
      type_cast_1232_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1232_inst_req_1;
      type_cast_1232_inst_ack_1<= rack(0);
      type_cast_1232_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1232_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1231_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv164_1233,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1249_inst_req_0;
      type_cast_1249_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1249_inst_req_1;
      type_cast_1249_inst_ack_1<= rack(0);
      type_cast_1249_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add144_1194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1249_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1256_inst_req_0;
      type_cast_1256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1256_inst_req_1;
      type_cast_1256_inst_ack_1<= rack(0);
      type_cast_1256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1256_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1258_inst_req_0;
      type_cast_1258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1258_inst_req_1;
      type_cast_1258_inst_ack_1<= rack(0);
      type_cast_1258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc161x_xix_x2_1221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1258_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1262_inst_req_0;
      type_cast_1262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1262_inst_req_1;
      type_cast_1262_inst_ack_1<= rack(0);
      type_cast_1262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1262_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1264_inst_req_0;
      type_cast_1264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1264_inst_req_1;
      type_cast_1264_inst_ack_1<= rack(0);
      type_cast_1264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1264_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_796_inst_req_0;
      type_cast_796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_796_inst_req_1;
      type_cast_796_inst_ack_1<= rack(0);
      type_cast_796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_800_inst_req_0;
      type_cast_800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_800_inst_req_1;
      type_cast_800_inst_ack_1<= rack(0);
      type_cast_800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_804_inst_req_0;
      type_cast_804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_804_inst_req_1;
      type_cast_804_inst_ack_1<= rack(0);
      type_cast_804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_805,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_808_inst_req_0;
      type_cast_808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_808_inst_req_1;
      type_cast_808_inst_ack_1<= rack(0);
      type_cast_808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_809,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_821_inst_req_0;
      type_cast_821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_821_inst_req_1;
      type_cast_821_inst_ack_1<= rack(0);
      type_cast_821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_822,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_831_inst
    process(sext185_828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext185_828(31 downto 0);
      type_cast_831_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_836_inst
    process(ASHR_i32_i32_835_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_835_wire(31 downto 0);
      conv82_837 <= tmp_var; -- 
    end process;
    type_cast_857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_857_inst_req_0;
      type_cast_857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_857_inst_req_1;
      type_cast_857_inst_ack_1<= rack(0);
      type_cast_857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_774,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_893_inst
    process(sext_890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_890(31 downto 0);
      type_cast_893_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_898_inst
    process(ASHR_i32_i32_897_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_897_wire(31 downto 0);
      conv100_899 <= tmp_var; -- 
    end process;
    type_cast_909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_909_inst_req_0;
      type_cast_909_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_909_inst_req_1;
      type_cast_909_inst_ack_1<= rack(0);
      type_cast_909_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_909_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_916_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_928_inst_req_0;
      type_cast_928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_928_inst_req_1;
      type_cast_928_inst_ack_1<= rack(0);
      type_cast_928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_927_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_929,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_932_inst
    process(conv42_929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv42_929(31 downto 0);
      type_cast_932_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_934_inst
    process(conv44_818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv44_818(31 downto 0);
      type_cast_934_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_945_inst
    process(conv42_929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv42_929(31 downto 0);
      type_cast_945_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_947_inst
    process(add_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_874(31 downto 0);
      type_cast_947_wire <= tmp_var; -- 
    end process;
    type_cast_965_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_965_inst_req_0;
      type_cast_965_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_965_inst_req_1;
      type_cast_965_inst_ack_1<= rack(0);
      type_cast_965_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_965_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_964_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_966,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_969_inst
    process(conv56_966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv56_966(31 downto 0);
      type_cast_969_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_971_inst
    process(conv44_818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv44_818(31 downto 0);
      type_cast_971_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_982_inst
    process(conv56_966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv56_966(31 downto 0);
      type_cast_982_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_984_inst
    process(add69_879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add69_879(31 downto 0);
      type_cast_984_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_1047_index_1_rename
    process(R_idxprom_1046_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1046_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1046_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1047_index_1_resize
    process(idxprom_1042) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1042;
      ov := iv(13 downto 0);
      R_idxprom_1046_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1047_root_address_inst
    process(array_obj_ref_1047_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1047_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1047_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1130_index_1_rename
    process(R_idxprom126_1129_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom126_1129_resized;
      ov(13 downto 0) := iv;
      R_idxprom126_1129_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1130_index_1_resize
    process(idxprom126_1125) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom126_1125;
      ov := iv(13 downto 0);
      R_idxprom126_1129_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1130_root_address_inst
    process(array_obj_ref_1130_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1130_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1130_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_index_1_rename
    process(R_idxprom131_1154_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom131_1154_resized;
      ov(13 downto 0) := iv;
      R_idxprom131_1154_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_index_1_resize
    process(idxprom131_1150) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom131_1150;
      ov := iv(13 downto 0);
      R_idxprom131_1154_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_root_address_inst
    process(array_obj_ref_1155_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1155_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1155_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1051_addr_0
    process(ptr_deref_1051_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1051_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1051_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1051_base_resize
    process(arrayidx_1049) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1049;
      ov := iv(13 downto 0);
      ptr_deref_1051_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1051_gather_scatter
    process(type_cast_1053_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1053_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1051_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1051_root_address_inst
    process(ptr_deref_1051_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1051_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1051_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1135_addr_0
    process(ptr_deref_1135_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1135_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1135_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1135_base_resize
    process(arrayidx127_1132) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx127_1132;
      ov := iv(13 downto 0);
      ptr_deref_1135_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1135_gather_scatter
    process(ptr_deref_1135_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1135_data_0;
      ov(63 downto 0) := iv;
      tmp128_1136 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1135_root_address_inst
    process(ptr_deref_1135_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1135_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1135_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1159_addr_0
    process(ptr_deref_1159_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1159_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1159_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1159_base_resize
    process(arrayidx132_1157) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx132_1157;
      ov := iv(13 downto 0);
      ptr_deref_1159_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1159_gather_scatter
    process(tmp128_1136) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp128_1136;
      ov(63 downto 0) := iv;
      ptr_deref_1159_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1159_root_address_inst
    process(ptr_deref_1159_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1159_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1159_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1182_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp139_1181;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1182_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1182_branch_req_0,
          ack0 => if_stmt_1182_branch_ack_0,
          ack1 => if_stmt_1182_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1239_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp172_1238;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1239_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1239_branch_req_0,
          ack0 => if_stmt_1239_branch_ack_0,
          ack1 => if_stmt_1239_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_955_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_954;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_955_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_955_branch_req_0,
          ack0 => if_stmt_955_branch_ack_0,
          ack1 => if_stmt_955_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_992_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond186_991;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_992_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_992_branch_req_0,
          ack0 => if_stmt_992_branch_ack_0,
          ack1 => if_stmt_992_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1193_inst
    process(kx_x1_902) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_902, type_cast_1192_wire_constant, tmp_var);
      add144_1194 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1201_inst
    process(jx_x1_917) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_917, type_cast_1200_wire_constant, tmp_var);
      inc_1202 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1220_inst
    process(inc161_1216, ix_x2_910) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc161_1216, ix_x2_910, tmp_var);
      inc161x_xix_x2_1221 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1022_inst
    process(mul85_1018, conv74_1003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul85_1018, conv74_1003, tmp_var);
      add80_1023 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1027_inst
    process(add80_1023, mul79_1013) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add80_1023, mul79_1013, tmp_var);
      add86_1028 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1085_inst
    process(mul106_1081, conv90_1061) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul106_1081, conv90_1061, tmp_var);
      add98_1086 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1090_inst
    process(add98_1086, mul97_1071) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add98_1086, mul97_1071, tmp_var);
      add107_1091 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1105_inst
    process(mul122_1101, conv90_1061) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul122_1101, conv90_1061, tmp_var);
      add117_1106 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1110_inst
    process(add117_1106, mul116_1096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add117_1106, mul116_1096, tmp_var);
      add123_1111 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1173_inst
    process(conv135_1168) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv135_1168, type_cast_1172_wire_constant, tmp_var);
      add136_1174 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_853_inst
    process(shl_849, div152_843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_849, div152_843, tmp_var);
      add155_854 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_868_inst
    process(shl_849, div167_864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_849, div167_864, tmp_var);
      add171_869 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_873_inst
    process(conv44_818, div167_864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv44_818, div167_864, tmp_var);
      add_874 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_878_inst
    process(conv44_818, div152_843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv44_818, div152_843, tmp_var);
      add69_879 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_953_inst
    process(cmpx_xnot_942, cmp52_949) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_942, cmp52_949, tmp_var);
      orx_xcond_954 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_990_inst
    process(cmp59x_xnot_979, cmp70_986) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp59x_xnot_979, cmp70_986, tmp_var);
      orx_xcond186_991 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1035_inst
    process(type_cast_1031_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1031_wire, type_cast_1034_wire_constant, tmp_var);
      ASHR_i32_i32_1035_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1118_inst
    process(type_cast_1114_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1114_wire, type_cast_1117_wire_constant, tmp_var);
      ASHR_i32_i32_1118_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1143_inst
    process(type_cast_1139_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1139_wire, type_cast_1142_wire_constant, tmp_var);
      ASHR_i32_i32_1143_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_835_inst
    process(type_cast_831_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_831_wire, type_cast_834_wire_constant, tmp_var);
      ASHR_i32_i32_835_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_897_inst
    process(type_cast_893_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_893_wire, type_cast_896_wire_constant, tmp_var);
      ASHR_i32_i32_897_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1211_inst
    process(conv149_1207, add155_854) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv149_1207, add155_854, tmp_var);
      cmp156_1212 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1237_inst
    process(conv164_1233, add171_869) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv164_1233, add171_869, tmp_var);
      cmp172_1238 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_842_inst
    process(conv29_801) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv29_801, type_cast_841_wire_constant, tmp_var);
      div152_843 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_863_inst
    process(conv166_858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv166_858, type_cast_862_wire_constant, tmp_var);
      div167_864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1012_inst
    process(conv78_1008, conv76_822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv78_1008, conv76_822, tmp_var);
      mul79_1013 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1017_inst
    process(conv42_929, conv82_837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_929, conv82_837, tmp_var);
      mul85_1018 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1070_inst
    process(sub_1066, conv27_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1066, conv27_797, tmp_var);
      mul97_1071 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1080_inst
    process(sub105_1076, conv100_899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub105_1076, conv100_899, tmp_var);
      mul106_1081 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1095_inst
    process(conv56_966, conv76_822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv56_966, conv76_822, tmp_var);
      mul116_1096 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1100_inst
    process(conv42_929, conv82_837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_929, conv82_837, tmp_var);
      mul122_1101 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_813_inst
    process(conv33_805, conv35_809) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_805, conv35_809, tmp_var);
      mul36_814 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_889_inst
    process(mul_885, conv27_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_885, conv27_797, tmp_var);
      sext_890 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_827_inst
    process(mul36_814) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul36_814, type_cast_826_wire_constant, tmp_var);
      sext185_828 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_848_inst
    process(conv44_818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_818, type_cast_847_wire_constant, tmp_var);
      shl_849 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_884_inst
    process(conv29_801) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_801, type_cast_883_wire_constant, tmp_var);
      mul_885 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1180_inst
    process(type_cast_1177_wire, type_cast_1179_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1177_wire, type_cast_1179_wire, tmp_var);
      cmp139_1181 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_935_inst
    process(type_cast_932_wire, type_cast_934_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_932_wire, type_cast_934_wire, tmp_var);
      cmp_936 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_948_inst
    process(type_cast_945_wire, type_cast_947_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_945_wire, type_cast_947_wire, tmp_var);
      cmp52_949 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_972_inst
    process(type_cast_969_wire, type_cast_971_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_969_wire, type_cast_971_wire, tmp_var);
      cmp59_973 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_985_inst
    process(type_cast_982_wire, type_cast_984_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_982_wire, type_cast_984_wire, tmp_var);
      cmp70_986 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1065_inst
    process(conv56_966, conv44_818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv56_966, conv44_818, tmp_var);
      sub_1066 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1075_inst
    process(conv42_929, conv44_818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv42_929, conv44_818, tmp_var);
      sub105_1076 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_941_inst
    process(cmp_936) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_936, type_cast_940_wire_constant, tmp_var);
      cmpx_xnot_942 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_978_inst
    process(cmp59_973) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp59_973, type_cast_977_wire_constant, tmp_var);
      cmp59x_xnot_979 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_1047_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1046_scaled;
      array_obj_ref_1047_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1047_index_offset_req_0;
      array_obj_ref_1047_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1047_index_offset_req_1;
      array_obj_ref_1047_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_1130_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom126_1129_scaled;
      array_obj_ref_1130_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1130_index_offset_req_0;
      array_obj_ref_1130_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1130_index_offset_req_1;
      array_obj_ref_1130_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_1155_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom131_1154_scaled;
      array_obj_ref_1155_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1155_index_offset_req_0;
      array_obj_ref_1155_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1155_index_offset_req_1;
      array_obj_ref_1155_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- unary operator type_cast_1001_inst
    process(kx_x1_902) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_902, tmp_var);
      type_cast_1001_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1006_inst
    process(jx_x1_917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_917, tmp_var);
      type_cast_1006_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1040_inst
    process(shr_1037) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1037, tmp_var);
      type_cast_1040_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1059_inst
    process(kx_x1_902) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_902, tmp_var);
      type_cast_1059_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1123_inst
    process(shr125_1120) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr125_1120, tmp_var);
      type_cast_1123_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1148_inst
    process(shr130_1145) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr130_1145, tmp_var);
      type_cast_1148_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1166_inst
    process(kx_x1_902) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_902, tmp_var);
      type_cast_1166_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1205_inst
    process(inc_1202) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1202, tmp_var);
      type_cast_1205_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1231_inst
    process(inc161x_xix_x2_1221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc161x_xix_x2_1221, tmp_var);
      type_cast_1231_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_927_inst
    process(ix_x2_910) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_910, tmp_var);
      type_cast_927_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_964_inst
    process(jx_x1_917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_917, tmp_var);
      type_cast_964_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1135_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1135_load_0_req_0;
      ptr_deref_1135_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1135_load_0_req_1;
      ptr_deref_1135_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1135_word_address_0;
      ptr_deref_1135_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1159_store_0 ptr_deref_1051_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1159_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1051_store_0_req_0;
      ptr_deref_1159_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1051_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1159_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1051_store_0_req_1;
      ptr_deref_1159_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1051_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1159_word_address_0 & ptr_deref_1051_word_address_0;
      data_in <= ptr_deref_1159_data_0 & ptr_deref_1051_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_starting_773_inst RPIPE_Block0_starting_776_inst RPIPE_Block0_starting_779_inst RPIPE_Block0_starting_782_inst RPIPE_Block0_starting_785_inst RPIPE_Block0_starting_788_inst RPIPE_Block0_starting_791_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block0_starting_773_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_starting_776_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_starting_779_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_starting_782_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_starting_785_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_starting_788_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_starting_791_inst_req_0;
      RPIPE_Block0_starting_773_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_starting_776_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_starting_779_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_starting_782_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_starting_785_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_starting_788_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_starting_791_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block0_starting_773_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_starting_776_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_starting_779_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_starting_782_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_starting_785_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_starting_788_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_starting_791_inst_req_1;
      RPIPE_Block0_starting_773_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_starting_776_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_starting_779_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_starting_782_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_starting_785_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_starting_788_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_starting_791_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call_774 <= data_out(55 downto 48);
      call1_777 <= data_out(47 downto 40);
      call2_780 <= data_out(39 downto 32);
      call3_783 <= data_out(31 downto 24);
      call4_786 <= data_out(23 downto 16);
      call5_789 <= data_out(15 downto 8);
      call6_792 <= data_out(7 downto 0);
      Block0_starting_read_0_gI: SplitGuardInterface generic map(name => "Block0_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block0_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_starting_pipe_read_req(0),
          oack => Block0_starting_pipe_read_ack(0),
          odata => Block0_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_complete_1269_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_complete_1269_inst_req_0;
      WPIPE_Block0_complete_1269_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_complete_1269_inst_req_1;
      WPIPE_Block0_complete_1269_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1271_wire_constant;
      Block0_complete_write_0_gI: SplitGuardInterface generic map(name => "Block0_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_complete_pipe_write_req(0),
          oack => Block0_complete_pipe_write_ack(0),
          odata => Block0_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_A_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_B is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block1_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_B;
architecture zeropad3D_B_arch of zeropad3D_B is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_B_CP_3564_start: Boolean;
  signal zeropad3D_B_CP_3564_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1334_inst_req_0 : boolean;
  signal array_obj_ref_1556_index_offset_req_0 : boolean;
  signal type_cast_1569_inst_ack_0 : boolean;
  signal type_cast_1550_inst_ack_1 : boolean;
  signal addr_of_1557_final_reg_ack_1 : boolean;
  signal type_cast_1658_inst_ack_0 : boolean;
  signal type_cast_1658_inst_req_0 : boolean;
  signal if_stmt_1464_branch_ack_1 : boolean;
  signal addr_of_1640_final_reg_req_1 : boolean;
  signal type_cast_1368_inst_ack_0 : boolean;
  signal ptr_deref_1644_load_0_ack_0 : boolean;
  signal array_obj_ref_1639_index_offset_req_1 : boolean;
  signal type_cast_1633_inst_ack_0 : boolean;
  signal addr_of_1640_final_reg_req_0 : boolean;
  signal addr_of_1640_final_reg_ack_0 : boolean;
  signal type_cast_1334_inst_ack_0 : boolean;
  signal type_cast_1633_inst_req_1 : boolean;
  signal type_cast_1633_inst_ack_1 : boolean;
  signal array_obj_ref_1639_index_offset_ack_1 : boolean;
  signal type_cast_1334_inst_req_1 : boolean;
  signal type_cast_1633_inst_req_0 : boolean;
  signal addr_of_1640_final_reg_ack_1 : boolean;
  signal type_cast_1338_inst_ack_0 : boolean;
  signal type_cast_1338_inst_req_0 : boolean;
  signal array_obj_ref_1639_index_offset_req_0 : boolean;
  signal type_cast_1569_inst_req_1 : boolean;
  signal ptr_deref_1560_store_0_ack_0 : boolean;
  signal type_cast_1511_inst_req_0 : boolean;
  signal ptr_deref_1644_load_0_req_0 : boolean;
  signal array_obj_ref_1639_index_offset_ack_0 : boolean;
  signal ptr_deref_1560_store_0_ack_1 : boolean;
  signal ptr_deref_1644_load_0_ack_1 : boolean;
  signal ptr_deref_1644_load_0_req_1 : boolean;
  signal type_cast_1511_inst_ack_0 : boolean;
  signal ptr_deref_1560_store_0_req_1 : boolean;
  signal type_cast_1334_inst_ack_1 : boolean;
  signal type_cast_1550_inst_req_1 : boolean;
  signal type_cast_1511_inst_req_1 : boolean;
  signal type_cast_1569_inst_ack_1 : boolean;
  signal type_cast_1437_inst_req_0 : boolean;
  signal if_stmt_1464_branch_ack_0 : boolean;
  signal type_cast_1511_inst_ack_1 : boolean;
  signal type_cast_1437_inst_ack_0 : boolean;
  signal ptr_deref_1560_store_0_req_0 : boolean;
  signal type_cast_1474_inst_req_1 : boolean;
  signal type_cast_1474_inst_req_0 : boolean;
  signal type_cast_1658_inst_req_1 : boolean;
  signal type_cast_1658_inst_ack_1 : boolean;
  signal addr_of_1557_final_reg_req_1 : boolean;
  signal type_cast_1368_inst_req_0 : boolean;
  signal type_cast_1368_inst_ack_1 : boolean;
  signal type_cast_1368_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1280_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1280_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1280_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1280_inst_ack_1 : boolean;
  signal addr_of_1557_final_reg_ack_0 : boolean;
  signal addr_of_1557_final_reg_req_0 : boolean;
  signal if_stmt_1464_branch_req_0 : boolean;
  signal RPIPE_Block1_starting_1283_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1283_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1283_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1283_inst_ack_1 : boolean;
  signal type_cast_1569_inst_req_0 : boolean;
  signal type_cast_1550_inst_ack_0 : boolean;
  signal type_cast_1550_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1286_inst_req_0 : boolean;
  signal if_stmt_1501_branch_ack_0 : boolean;
  signal RPIPE_Block1_starting_1286_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1286_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1286_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1289_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1289_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1289_inst_req_1 : boolean;
  signal if_stmt_1501_branch_ack_1 : boolean;
  signal RPIPE_Block1_starting_1289_inst_ack_1 : boolean;
  signal type_cast_1516_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1292_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1292_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1292_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1292_inst_ack_1 : boolean;
  signal array_obj_ref_1556_index_offset_ack_1 : boolean;
  signal type_cast_1516_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1295_inst_req_0 : boolean;
  signal if_stmt_1501_branch_req_0 : boolean;
  signal RPIPE_Block1_starting_1295_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1295_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1295_inst_ack_1 : boolean;
  signal array_obj_ref_1556_index_offset_req_1 : boolean;
  signal type_cast_1516_inst_ack_0 : boolean;
  signal type_cast_1516_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1298_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1298_inst_ack_0 : boolean;
  signal type_cast_1338_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1298_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1298_inst_ack_1 : boolean;
  signal array_obj_ref_1556_index_offset_ack_0 : boolean;
  signal type_cast_1303_inst_req_0 : boolean;
  signal type_cast_1303_inst_ack_0 : boolean;
  signal type_cast_1474_inst_ack_0 : boolean;
  signal type_cast_1303_inst_req_1 : boolean;
  signal type_cast_1474_inst_ack_1 : boolean;
  signal type_cast_1303_inst_ack_1 : boolean;
  signal type_cast_1338_inst_req_1 : boolean;
  signal type_cast_1437_inst_ack_1 : boolean;
  signal type_cast_1437_inst_req_1 : boolean;
  signal type_cast_1313_inst_req_0 : boolean;
  signal type_cast_1313_inst_ack_0 : boolean;
  signal type_cast_1313_inst_req_1 : boolean;
  signal type_cast_1313_inst_ack_1 : boolean;
  signal type_cast_1317_inst_req_0 : boolean;
  signal type_cast_1317_inst_ack_0 : boolean;
  signal type_cast_1317_inst_req_1 : boolean;
  signal type_cast_1317_inst_ack_1 : boolean;
  signal type_cast_1321_inst_req_0 : boolean;
  signal type_cast_1321_inst_ack_0 : boolean;
  signal type_cast_1321_inst_req_1 : boolean;
  signal type_cast_1321_inst_ack_1 : boolean;
  signal type_cast_1325_inst_req_0 : boolean;
  signal type_cast_1325_inst_ack_0 : boolean;
  signal type_cast_1325_inst_req_1 : boolean;
  signal type_cast_1325_inst_ack_1 : boolean;
  signal array_obj_ref_1664_index_offset_req_0 : boolean;
  signal array_obj_ref_1664_index_offset_ack_0 : boolean;
  signal array_obj_ref_1664_index_offset_req_1 : boolean;
  signal array_obj_ref_1664_index_offset_ack_1 : boolean;
  signal addr_of_1665_final_reg_req_0 : boolean;
  signal addr_of_1665_final_reg_ack_0 : boolean;
  signal addr_of_1665_final_reg_req_1 : boolean;
  signal addr_of_1665_final_reg_ack_1 : boolean;
  signal ptr_deref_1668_store_0_req_0 : boolean;
  signal ptr_deref_1668_store_0_ack_0 : boolean;
  signal ptr_deref_1668_store_0_req_1 : boolean;
  signal ptr_deref_1668_store_0_ack_1 : boolean;
  signal type_cast_1676_inst_req_0 : boolean;
  signal type_cast_1676_inst_ack_0 : boolean;
  signal type_cast_1676_inst_req_1 : boolean;
  signal type_cast_1676_inst_ack_1 : boolean;
  signal if_stmt_1691_branch_req_0 : boolean;
  signal if_stmt_1691_branch_ack_1 : boolean;
  signal if_stmt_1691_branch_ack_0 : boolean;
  signal type_cast_1715_inst_req_0 : boolean;
  signal type_cast_1715_inst_ack_0 : boolean;
  signal type_cast_1715_inst_req_1 : boolean;
  signal type_cast_1715_inst_ack_1 : boolean;
  signal type_cast_1724_inst_req_0 : boolean;
  signal type_cast_1724_inst_ack_0 : boolean;
  signal type_cast_1724_inst_req_1 : boolean;
  signal type_cast_1724_inst_ack_1 : boolean;
  signal type_cast_1740_inst_req_0 : boolean;
  signal type_cast_1740_inst_ack_0 : boolean;
  signal type_cast_1740_inst_req_1 : boolean;
  signal type_cast_1740_inst_ack_1 : boolean;
  signal if_stmt_1747_branch_req_0 : boolean;
  signal if_stmt_1747_branch_ack_1 : boolean;
  signal if_stmt_1747_branch_ack_0 : boolean;
  signal WPIPE_Block1_complete_1777_inst_req_0 : boolean;
  signal WPIPE_Block1_complete_1777_inst_ack_0 : boolean;
  signal WPIPE_Block1_complete_1777_inst_req_1 : boolean;
  signal WPIPE_Block1_complete_1777_inst_ack_1 : boolean;
  signal phi_stmt_1413_req_0 : boolean;
  signal phi_stmt_1420_req_0 : boolean;
  signal type_cast_1430_inst_req_0 : boolean;
  signal type_cast_1430_inst_ack_0 : boolean;
  signal type_cast_1430_inst_req_1 : boolean;
  signal type_cast_1430_inst_ack_1 : boolean;
  signal phi_stmt_1427_req_0 : boolean;
  signal type_cast_1419_inst_req_0 : boolean;
  signal type_cast_1419_inst_ack_0 : boolean;
  signal type_cast_1419_inst_req_1 : boolean;
  signal type_cast_1419_inst_ack_1 : boolean;
  signal phi_stmt_1413_req_1 : boolean;
  signal type_cast_1426_inst_req_0 : boolean;
  signal type_cast_1426_inst_ack_0 : boolean;
  signal type_cast_1426_inst_req_1 : boolean;
  signal type_cast_1426_inst_ack_1 : boolean;
  signal phi_stmt_1420_req_1 : boolean;
  signal type_cast_1432_inst_req_0 : boolean;
  signal type_cast_1432_inst_ack_0 : boolean;
  signal type_cast_1432_inst_req_1 : boolean;
  signal type_cast_1432_inst_ack_1 : boolean;
  signal phi_stmt_1427_req_1 : boolean;
  signal phi_stmt_1413_ack_0 : boolean;
  signal phi_stmt_1420_ack_0 : boolean;
  signal phi_stmt_1427_ack_0 : boolean;
  signal type_cast_1766_inst_req_0 : boolean;
  signal type_cast_1766_inst_ack_0 : boolean;
  signal type_cast_1766_inst_req_1 : boolean;
  signal type_cast_1766_inst_ack_1 : boolean;
  signal phi_stmt_1761_req_1 : boolean;
  signal type_cast_1772_inst_req_0 : boolean;
  signal type_cast_1772_inst_ack_0 : boolean;
  signal type_cast_1772_inst_req_1 : boolean;
  signal type_cast_1772_inst_ack_1 : boolean;
  signal phi_stmt_1767_req_1 : boolean;
  signal phi_stmt_1754_req_1 : boolean;
  signal type_cast_1764_inst_req_0 : boolean;
  signal type_cast_1764_inst_ack_0 : boolean;
  signal type_cast_1764_inst_req_1 : boolean;
  signal type_cast_1764_inst_ack_1 : boolean;
  signal phi_stmt_1761_req_0 : boolean;
  signal type_cast_1770_inst_req_0 : boolean;
  signal type_cast_1770_inst_ack_0 : boolean;
  signal type_cast_1770_inst_req_1 : boolean;
  signal type_cast_1770_inst_ack_1 : boolean;
  signal phi_stmt_1767_req_0 : boolean;
  signal type_cast_1757_inst_req_0 : boolean;
  signal type_cast_1757_inst_ack_0 : boolean;
  signal type_cast_1757_inst_req_1 : boolean;
  signal type_cast_1757_inst_ack_1 : boolean;
  signal phi_stmt_1754_req_0 : boolean;
  signal phi_stmt_1754_ack_0 : boolean;
  signal phi_stmt_1761_ack_0 : boolean;
  signal phi_stmt_1767_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_B_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_B_CP_3564_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_B_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_B_CP_3564_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_B_CP_3564_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_B_CP_3564_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_B_CP_3564: Block -- control-path 
    signal zeropad3D_B_CP_3564_elements: BooleanArray(134 downto 0);
    -- 
  begin -- 
    zeropad3D_B_CP_3564_elements(0) <= zeropad3D_B_CP_3564_start;
    zeropad3D_B_CP_3564_symbol <= zeropad3D_B_CP_3564_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1278/$entry
      -- CP-element group 0: 	 branch_block_stmt_1278/branch_block_stmt_1278__entry__
      -- CP-element group 0: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299__entry__
      -- CP-element group 0: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/$entry
      -- CP-element group 0: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Sample/rr
      -- 
    rr_3630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(0), ack => RPIPE_Block1_starting_1280_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	134 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	102 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_1278/merge_stmt_1753__exit__
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Update/cr
      -- 
    rr_4466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(1), ack => type_cast_1419_inst_req_0); -- 
    cr_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(1), ack => type_cast_1419_inst_req_1); -- 
    rr_4489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(1), ack => type_cast_1426_inst_req_0); -- 
    cr_4494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(1), ack => type_cast_1426_inst_req_1); -- 
    rr_4512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(1), ack => type_cast_1432_inst_req_0); -- 
    cr_4517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(1), ack => type_cast_1432_inst_req_1); -- 
    zeropad3D_B_CP_3564_elements(1) <= zeropad3D_B_CP_3564_elements(134);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Update/cr
      -- 
    ra_3631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1280_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(2)); -- 
    cr_3635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(2), ack => RPIPE_Block1_starting_1280_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1280_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Sample/rr
      -- 
    ca_3636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1280_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(3)); -- 
    rr_3644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(3), ack => RPIPE_Block1_starting_1283_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Update/cr
      -- 
    ra_3645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1283_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(4)); -- 
    cr_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(4), ack => RPIPE_Block1_starting_1283_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1283_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Sample/rr
      -- 
    ca_3650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1283_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(5)); -- 
    rr_3658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(5), ack => RPIPE_Block1_starting_1286_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Update/cr
      -- 
    ra_3659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1286_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(6)); -- 
    cr_3663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(6), ack => RPIPE_Block1_starting_1286_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1286_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Sample/rr
      -- 
    ca_3664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1286_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(7)); -- 
    rr_3672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(7), ack => RPIPE_Block1_starting_1289_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Update/cr
      -- 
    ra_3673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1289_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(8)); -- 
    cr_3677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(8), ack => RPIPE_Block1_starting_1289_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1289_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Sample/rr
      -- 
    ca_3678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1289_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(9)); -- 
    rr_3686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(9), ack => RPIPE_Block1_starting_1292_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Update/cr
      -- 
    ra_3687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1292_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(10)); -- 
    cr_3691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(10), ack => RPIPE_Block1_starting_1292_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1292_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Sample/rr
      -- 
    ca_3692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1292_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(11)); -- 
    rr_3700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(11), ack => RPIPE_Block1_starting_1295_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Update/cr
      -- 
    ra_3701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1295_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(12)); -- 
    cr_3705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(12), ack => RPIPE_Block1_starting_1295_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1295_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Sample/rr
      -- 
    ca_3706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1295_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(13)); -- 
    rr_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(13), ack => RPIPE_Block1_starting_1298_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Update/cr
      -- 
    ra_3715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1298_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(14)); -- 
    cr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(14), ack => RPIPE_Block1_starting_1298_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15:  members (55) 
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299__exit__
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410__entry__
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/$exit
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1281_to_assign_stmt_1299/RPIPE_Block1_starting_1298_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_update_start_
      -- 
    ca_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1298_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(15)); -- 
    rr_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1334_inst_req_0); -- 
    cr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1334_inst_req_1); -- 
    rr_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1338_inst_req_0); -- 
    rr_3829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1368_inst_req_0); -- 
    cr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1368_inst_req_1); -- 
    rr_3731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1303_inst_req_0); -- 
    cr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1303_inst_req_1); -- 
    cr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1338_inst_req_1); -- 
    rr_3745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1313_inst_req_0); -- 
    cr_3750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1313_inst_req_1); -- 
    rr_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1317_inst_req_0); -- 
    cr_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1317_inst_req_1); -- 
    rr_3773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1321_inst_req_0); -- 
    cr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1321_inst_req_1); -- 
    rr_3787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1325_inst_req_0); -- 
    cr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(15), ack => type_cast_1325_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Sample/ra
      -- 
    ra_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1303_Update/ca
      -- 
    ca_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Sample/ra
      -- 
    ra_3746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1313_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1313_Update/ca
      -- 
    ca_3751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1313_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Sample/ra
      -- 
    ra_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1317_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1317_Update/ca
      -- 
    ca_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1317_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Sample/ra
      -- 
    ra_3774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1321_Update/ca
      -- 
    ca_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Sample/ra
      -- 
    ra_3788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1325_Update/ca
      -- 
    ca_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_sample_completed_
      -- 
    ra_3802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1334_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1334_update_completed_
      -- 
    ca_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1334_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Sample/$exit
      -- 
    ra_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1338_Update/$exit
      -- 
    ca_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_sample_completed_
      -- 
    ra_3830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/type_cast_1368_update_completed_
      -- 
    ca_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	21 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	25 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: 	90 
    -- CP-element group 32: 	91 
    -- CP-element group 32: 	92 
    -- CP-element group 32:  members (16) 
      -- CP-element group 32: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410__exit__
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody
      -- CP-element group 32: 	 branch_block_stmt_1278/assign_stmt_1304_to_assign_stmt_1410/$exit
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1413/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1420/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/cr
      -- 
    rr_4440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(32), ack => type_cast_1430_inst_req_0); -- 
    cr_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(32), ack => type_cast_1430_inst_req_1); -- 
    zeropad3D_B_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(17) & zeropad3D_B_CP_3564_elements(19) & zeropad3D_B_CP_3564_elements(21) & zeropad3D_B_CP_3564_elements(23) & zeropad3D_B_CP_3564_elements(25) & zeropad3D_B_CP_3564_elements(27) & zeropad3D_B_CP_3564_elements(29) & zeropad3D_B_CP_3564_elements(31);
      gj_zeropad3D_B_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	109 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_sample_completed_
      -- 
    ra_3847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	109 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (13) 
      -- CP-element group 34: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464_else_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463__exit__
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464__entry__
      -- CP-element group 34: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/$exit
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464_eval_test/branch_req
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_1278/if_stmt_1464_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1278/R_orx_xcond_1465_place
      -- 
    ca_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(34)); -- 
    branch_req_3860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(34), ack => if_stmt_1464_branch_req_0); -- 
    -- CP-element group 35:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (18) 
      -- CP-element group 35: 	 branch_block_stmt_1278/if_stmt_1464_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/$entry
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1278/if_stmt_1464_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_1278/merge_stmt_1470__exit__
      -- CP-element group 35: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500__entry__
      -- CP-element group 35: 	 branch_block_stmt_1278/whilex_xbody_lorx_xlhsx_xfalse60
      -- CP-element group 35: 	 branch_block_stmt_1278/whilex_xbody_lorx_xlhsx_xfalse60_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_1278/whilex_xbody_lorx_xlhsx_xfalse60_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_1278/merge_stmt_1470_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_1278/merge_stmt_1470_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_1278/merge_stmt_1470_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_1278/merge_stmt_1470_PhiAck/dummy
      -- 
    if_choice_transition_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1464_branch_ack_1, ack => zeropad3D_B_CP_3564_elements(35)); -- 
    cr_3887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(35), ack => type_cast_1474_inst_req_1); -- 
    rr_3882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(35), ack => type_cast_1474_inst_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	110 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1278/if_stmt_1464_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_1278/if_stmt_1464_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_1278/whilex_xbody_ifx_xthen
      -- CP-element group 36: 	 branch_block_stmt_1278/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1278/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1464_branch_ack_0, ack => zeropad3D_B_CP_3564_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Sample/ra
      -- 
    ra_3883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1474_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (13) 
      -- CP-element group 38: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/$exit
      -- CP-element group 38: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500__exit__
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501__entry__
      -- CP-element group 38: 	 branch_block_stmt_1278/R_orx_xcond190_1502_place
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501_else_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501_if_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501_eval_test/branch_req
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_1278/if_stmt_1501_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1278/assign_stmt_1475_to_assign_stmt_1500/type_cast_1474_Update/ca
      -- 
    ca_3888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1474_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(38)); -- 
    branch_req_3896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(38), ack => if_stmt_1501_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/merge_stmt_1565__exit__
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670__entry__
      -- CP-element group 39: 	 branch_block_stmt_1278/lorx_xlhsx_xfalse60_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/if_stmt_1501_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_1278/if_stmt_1501_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1278/lorx_xlhsx_xfalse60_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/lorx_xlhsx_xfalse60_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_1278/merge_stmt_1565_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_1278/merge_stmt_1565_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_1278/merge_stmt_1565_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_1278/merge_stmt_1565_PhiAck/dummy
      -- 
    if_choice_transition_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1501_branch_ack_1, ack => zeropad3D_B_CP_3564_elements(39)); -- 
    req_4124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => addr_of_1640_final_reg_req_1); -- 
    req_4109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => array_obj_ref_1639_index_offset_req_1); -- 
    cr_4078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => type_cast_1633_inst_req_1); -- 
    cr_4064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => type_cast_1569_inst_req_1); -- 
    cr_4169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => ptr_deref_1644_load_0_req_1); -- 
    cr_4188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => type_cast_1658_inst_req_1); -- 
    rr_4059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => type_cast_1569_inst_req_0); -- 
    req_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => array_obj_ref_1664_index_offset_req_1); -- 
    req_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => addr_of_1665_final_reg_req_1); -- 
    cr_4284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(39), ack => ptr_deref_1668_store_0_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	110 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1278/lorx_xlhsx_xfalse60_ifx_xthen
      -- CP-element group 40: 	 branch_block_stmt_1278/if_stmt_1501_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_1278/if_stmt_1501_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_1278/lorx_xlhsx_xfalse60_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_1278/lorx_xlhsx_xfalse60_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1501_branch_ack_0, ack => zeropad3D_B_CP_3564_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	110 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_sample_completed_
      -- 
    ra_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	110 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_update_completed_
      -- 
    ca_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	110 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_sample_completed_
      -- 
    ra_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1516_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Update/$exit
      -- 
    ca_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1516_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_sample_start_
      -- 
    rr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(45), ack => type_cast_1550_inst_req_0); -- 
    zeropad3D_B_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(44) & zeropad3D_B_CP_3564_elements(42);
      gj_zeropad3D_B_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_sample_completed_
      -- 
    ra_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	110 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_index_computed_1
      -- 
    ca_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(47)); -- 
    req_3977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(47), ack => array_obj_ref_1556_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Sample/ack
      -- 
    ack_3978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1556_index_offset_ack_0, ack => zeropad3D_B_CP_3564_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	110 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_request/req
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Update/$exit
      -- 
    ack_3983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1556_index_offset_ack_1, ack => zeropad3D_B_CP_3564_elements(49)); -- 
    req_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(49), ack => addr_of_1557_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_request/ack
      -- CP-element group 50: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_request/$exit
      -- 
    ack_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1557_final_reg_ack_0, ack => zeropad3D_B_CP_3564_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	110 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/ptr_deref_1560_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/word_access_start/word_0/rr
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/ptr_deref_1560_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/ptr_deref_1560_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/ptr_deref_1560_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_word_addrgen/$entry
      -- 
    ack_3998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1557_final_reg_ack_1, ack => zeropad3D_B_CP_3564_elements(51)); -- 
    rr_4036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(51), ack => ptr_deref_1560_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/word_access_start/word_0/ra
      -- CP-element group 52: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Sample/$exit
      -- 
    ra_4037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1560_store_0_ack_0, ack => zeropad3D_B_CP_3564_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	110 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_update_completed_
      -- 
    ca_4048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1560_store_0_ack_1, ack => zeropad3D_B_CP_3564_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	48 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	111 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563__exit__
      -- CP-element group 54: 	 branch_block_stmt_1278/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/$exit
      -- CP-element group 54: 	 branch_block_stmt_1278/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1278/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(48) & zeropad3D_B_CP_3564_elements(53);
      gj_zeropad3D_B_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Sample/$exit
      -- 
    ra_4060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1569_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1569_update_completed_
      -- 
    ca_4065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1569_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(56)); -- 
    rr_4073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(56), ack => type_cast_1633_inst_req_0); -- 
    rr_4183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(56), ack => type_cast_1658_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_sample_completed_
      -- 
    ra_4074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1633_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1633_update_completed_
      -- 
    ca_4079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1633_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(58)); -- 
    req_4104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(58), ack => array_obj_ref_1639_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_sample_complete
      -- 
    ack_4105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1639_index_offset_ack_0, ack => zeropad3D_B_CP_3564_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_request/req
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1639_base_plus_offset/sum_rename_ack
      -- 
    ack_4110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1639_index_offset_ack_1, ack => zeropad3D_B_CP_3564_elements(60)); -- 
    req_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(60), ack => addr_of_1640_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_request/ack
      -- CP-element group 61: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_request/$exit
      -- 
    ack_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1640_final_reg_ack_0, ack => zeropad3D_B_CP_3564_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/word_access_start/word_0/rr
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1640_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_base_address_resized
      -- 
    ack_4125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1640_final_reg_ack_1, ack => zeropad3D_B_CP_3564_elements(62)); -- 
    rr_4158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(62), ack => ptr_deref_1644_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/word_access_start/word_0/ra
      -- CP-element group 63: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Sample/word_access_start/word_0/$exit
      -- 
    ra_4159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1644_load_0_ack_0, ack => zeropad3D_B_CP_3564_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/ptr_deref_1644_Merge/merge_ack
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/ptr_deref_1644_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/ptr_deref_1644_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1644_Update/ptr_deref_1644_Merge/$entry
      -- 
    ca_4170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1644_load_0_ack_1, ack => zeropad3D_B_CP_3564_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_sample_completed_
      -- 
    ra_4184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/type_cast_1658_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_computed_1
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Sample/req
      -- 
    ca_4189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(66)); -- 
    req_4214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(66), ack => array_obj_ref_1664_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Sample/ack
      -- 
    ack_4215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1664_index_offset_ack_0, ack => zeropad3D_B_CP_3564_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/array_obj_ref_1664_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_request/req
      -- 
    ack_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1664_index_offset_ack_1, ack => zeropad3D_B_CP_3564_elements(68)); -- 
    req_4229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(68), ack => addr_of_1665_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_request/ack
      -- 
    ack_4230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1665_final_reg_ack_0, ack => zeropad3D_B_CP_3564_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/addr_of_1665_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_word_addrgen/root_register_ack
      -- 
    ack_4235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1665_final_reg_ack_1, ack => zeropad3D_B_CP_3564_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/ptr_deref_1668_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/ptr_deref_1668_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/ptr_deref_1668_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/ptr_deref_1668_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/word_access_start/word_0/rr
      -- 
    rr_4273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(71), ack => ptr_deref_1668_store_0_req_0); -- 
    zeropad3D_B_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(64) & zeropad3D_B_CP_3564_elements(70);
      gj_zeropad3D_B_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Sample/word_access_start/word_0/ra
      -- 
    ra_4274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1668_store_0_ack_0, ack => zeropad3D_B_CP_3564_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/ptr_deref_1668_Update/word_access_complete/word_0/ca
      -- 
    ca_4285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1668_store_0_ack_1, ack => zeropad3D_B_CP_3564_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	111 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670/$exit
      -- CP-element group 74: 	 branch_block_stmt_1278/assign_stmt_1570_to_assign_stmt_1670__exit__
      -- CP-element group 74: 	 branch_block_stmt_1278/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_1278/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_1278/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(59) & zeropad3D_B_CP_3564_elements(67) & zeropad3D_B_CP_3564_elements(73);
      gj_zeropad3D_B_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	111 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Sample/ra
      -- 
    ra_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	111 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_1278/R_cmp144_1692_place
      -- CP-element group 76: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690__exit__
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691__entry__
      -- CP-element group 76: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/$exit
      -- CP-element group 76: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1278/if_stmt_1691_else_link/$entry
      -- 
    ca_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(76)); -- 
    branch_req_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(76), ack => if_stmt_1691_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	127 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xend_ifx_xthen146
      -- CP-element group 77: 	 branch_block_stmt_1278/merge_stmt_1697__exit__
      -- CP-element group 77: 	 branch_block_stmt_1278/assign_stmt_1703__entry__
      -- CP-element group 77: 	 branch_block_stmt_1278/assign_stmt_1703__exit__
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184
      -- CP-element group 77: 	 branch_block_stmt_1278/if_stmt_1691_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_1278/if_stmt_1691_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_1278/assign_stmt_1703/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/assign_stmt_1703/$exit
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xend_ifx_xthen146_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xend_ifx_xthen146_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_1278/merge_stmt_1697_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_1278/merge_stmt_1697_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/merge_stmt_1697_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_1278/merge_stmt_1697_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1691_branch_ack_1, ack => zeropad3D_B_CP_3564_elements(77)); -- 
    rr_4672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(77), ack => type_cast_1764_inst_req_0); -- 
    cr_4677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(77), ack => type_cast_1764_inst_req_1); -- 
    rr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(77), ack => type_cast_1770_inst_req_0); -- 
    cr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(77), ack => type_cast_1770_inst_req_1); -- 
    rr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(77), ack => type_cast_1757_inst_req_0); -- 
    cr_4723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(77), ack => type_cast_1757_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (24) 
      -- CP-element group 78: 	 branch_block_stmt_1278/ifx_xend_ifx_xelse151
      -- CP-element group 78: 	 branch_block_stmt_1278/merge_stmt_1705__exit__
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746__entry__
      -- CP-element group 78: 	 branch_block_stmt_1278/if_stmt_1691_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_1278/if_stmt_1691_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1278/ifx_xend_ifx_xelse151_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/ifx_xend_ifx_xelse151_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1278/merge_stmt_1705_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1278/merge_stmt_1705_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1278/merge_stmt_1705_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1278/merge_stmt_1705_PhiAck/dummy
      -- 
    else_choice_transition_4319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1691_branch_ack_0, ack => zeropad3D_B_CP_3564_elements(78)); -- 
    rr_4335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(78), ack => type_cast_1715_inst_req_0); -- 
    cr_4340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(78), ack => type_cast_1715_inst_req_1); -- 
    cr_4354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(78), ack => type_cast_1724_inst_req_1); -- 
    cr_4368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(78), ack => type_cast_1740_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Sample/ra
      -- 
    ra_4336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1715_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1715_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Sample/rr
      -- 
    ca_4341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1715_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(80)); -- 
    rr_4349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(80), ack => type_cast_1724_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Sample/ra
      -- 
    ra_4350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1724_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Sample/rr
      -- 
    ca_4355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(82)); -- 
    rr_4363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(82), ack => type_cast_1740_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Sample/ra
      -- 
    ra_4364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1740_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(83)); -- 
    -- CP-element group 84:  branch  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (13) 
      -- CP-element group 84: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746__exit__
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747__entry__
      -- CP-element group 84: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/$exit
      -- CP-element group 84: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1278/assign_stmt_1711_to_assign_stmt_1746/type_cast_1740_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_1278/R_cmp176_1748_place
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1278/if_stmt_1747_else_link/$entry
      -- 
    ca_4369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1740_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(84)); -- 
    branch_req_4377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(84), ack => if_stmt_1747_branch_req_0); -- 
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_1278/merge_stmt_1775__exit__
      -- CP-element group 85: 	 branch_block_stmt_1278/assign_stmt_1780__entry__
      -- CP-element group 85: 	 branch_block_stmt_1278/if_stmt_1747_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_1278/if_stmt_1747_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_1278/ifx_xelse151_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_1278/assign_stmt_1780/$entry
      -- CP-element group 85: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_1278/ifx_xelse151_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_1278/ifx_xelse151_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1278/merge_stmt_1775_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1278/merge_stmt_1775_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_1278/merge_stmt_1775_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_1278/merge_stmt_1775_PhiAck/dummy
      -- 
    if_choice_transition_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1747_branch_ack_1, ack => zeropad3D_B_CP_3564_elements(85)); -- 
    req_4399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(85), ack => WPIPE_Block1_complete_1777_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	115 
    -- CP-element group 86: 	116 
    -- CP-element group 86: 	118 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_1278/if_stmt_1747_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_1278/if_stmt_1747_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1754/$entry
      -- CP-element group 86: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$entry
      -- 
    else_choice_transition_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1747_branch_ack_0, ack => zeropad3D_B_CP_3564_elements(86)); -- 
    rr_4615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(86), ack => type_cast_1766_inst_req_0); -- 
    cr_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(86), ack => type_cast_1766_inst_req_1); -- 
    rr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(86), ack => type_cast_1772_inst_req_0); -- 
    cr_4643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(86), ack => type_cast_1772_inst_req_1); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Update/req
      -- 
    ack_4400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_complete_1777_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(87)); -- 
    req_4404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(87), ack => WPIPE_Block1_complete_1777_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_1278/$exit
      -- CP-element group 88: 	 branch_block_stmt_1278/branch_block_stmt_1278__exit__
      -- CP-element group 88: 	 branch_block_stmt_1278/assign_stmt_1780__exit__
      -- CP-element group 88: 	 branch_block_stmt_1278/return__
      -- CP-element group 88: 	 branch_block_stmt_1278/merge_stmt_1782__exit__
      -- CP-element group 88: 	 branch_block_stmt_1278/assign_stmt_1780/$exit
      -- CP-element group 88: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1278/assign_stmt_1780/WPIPE_Block1_complete_1777_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1278/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_1278/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_1278/merge_stmt_1782_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1278/merge_stmt_1782_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_1278/merge_stmt_1782_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1278/merge_stmt_1782_PhiAck/dummy
      -- 
    ack_4405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_complete_1777_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(88)); -- 
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	94 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1413/$exit
      -- CP-element group 89: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1417_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_req
      -- 
    phi_stmt_1413_req_4416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1413_req_4416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(89), ack => phi_stmt_1413_req_0); -- 
    -- Element group zeropad3D_B_CP_3564_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_3564_elements(32), ack => zeropad3D_B_CP_3564_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	32 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1420/$exit
      -- CP-element group 90: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1424_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_req
      -- 
    phi_stmt_1420_req_4424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1420_req_4424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(90), ack => phi_stmt_1420_req_0); -- 
    -- Element group zeropad3D_B_CP_3564_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_3564_elements(32), ack => zeropad3D_B_CP_3564_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/ra
      -- 
    ra_4441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	32 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/ca
      -- 
    ca_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/$exit
      -- CP-element group 93: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/$exit
      -- CP-element group 93: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_req
      -- 
    phi_stmt_1427_req_4447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1427_req_4447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(93), ack => phi_stmt_1427_req_0); -- 
    zeropad3D_B_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(91) & zeropad3D_B_CP_3564_elements(92);
      gj_zeropad3D_B_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	105 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1278/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(89) & zeropad3D_B_CP_3564_elements(90) & zeropad3D_B_CP_3564_elements(93);
      gj_zeropad3D_B_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Sample/ra
      -- 
    ra_4467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1419_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/Update/ca
      -- 
    ca_4472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1419_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/$exit
      -- CP-element group 97: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/$exit
      -- CP-element group 97: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_sources/type_cast_1419/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1413/phi_stmt_1413_req
      -- 
    phi_stmt_1413_req_4473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1413_req_4473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(97), ack => phi_stmt_1413_req_1); -- 
    zeropad3D_B_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(95) & zeropad3D_B_CP_3564_elements(96);
      gj_zeropad3D_B_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Sample/ra
      -- 
    ra_4490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/Update/ca
      -- 
    ca_4495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/$exit
      -- CP-element group 100: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/$exit
      -- CP-element group 100: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_sources/type_cast_1426/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1420/phi_stmt_1420_req
      -- 
    phi_stmt_1420_req_4496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1420_req_4496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(100), ack => phi_stmt_1420_req_1); -- 
    zeropad3D_B_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(98) & zeropad3D_B_CP_3564_elements(99);
      gj_zeropad3D_B_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Sample/ra
      -- 
    ra_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1432_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/Update/ca
      -- 
    ca_4518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1432_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/$exit
      -- CP-element group 103: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/$exit
      -- CP-element group 103: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1432/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1427/phi_stmt_1427_req
      -- 
    phi_stmt_1427_req_4519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1427_req_4519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(103), ack => phi_stmt_1427_req_1); -- 
    zeropad3D_B_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(101) & zeropad3D_B_CP_3564_elements(102);
      gj_zeropad3D_B_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1278/ifx_xend184_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(97) & zeropad3D_B_CP_3564_elements(100) & zeropad3D_B_CP_3564_elements(103);
      gj_zeropad3D_B_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  merge  fork  transition  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	94 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1278/merge_stmt_1412_PhiReqMerge
      -- CP-element group 105: 	 branch_block_stmt_1278/merge_stmt_1412_PhiAck/$entry
      -- 
    zeropad3D_B_CP_3564_elements(105) <= OrReduce(zeropad3D_B_CP_3564_elements(94) & zeropad3D_B_CP_3564_elements(104));
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1278/merge_stmt_1412_PhiAck/phi_stmt_1413_ack
      -- 
    phi_stmt_1413_ack_4524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1413_ack_0, ack => zeropad3D_B_CP_3564_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1278/merge_stmt_1412_PhiAck/phi_stmt_1420_ack
      -- 
    phi_stmt_1420_ack_4525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1420_ack_0, ack => zeropad3D_B_CP_3564_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1278/merge_stmt_1412_PhiAck/phi_stmt_1427_ack
      -- 
    phi_stmt_1427_ack_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1427_ack_0, ack => zeropad3D_B_CP_3564_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	33 
    -- CP-element group 109: 	34 
    -- CP-element group 109:  members (10) 
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1278/merge_stmt_1412__exit__
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463__entry__
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/$entry
      -- CP-element group 109: 	 branch_block_stmt_1278/assign_stmt_1438_to_assign_stmt_1463/type_cast_1437_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_1278/merge_stmt_1412_PhiAck/$exit
      -- 
    rr_3846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(109), ack => type_cast_1437_inst_req_0); -- 
    cr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(109), ack => type_cast_1437_inst_req_1); -- 
    zeropad3D_B_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(106) & zeropad3D_B_CP_3564_elements(107) & zeropad3D_B_CP_3564_elements(108);
      gj_zeropad3D_B_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  merge  fork  transition  place  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	36 
    -- CP-element group 110: 	40 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	53 
    -- CP-element group 110: 	44 
    -- CP-element group 110: 	51 
    -- CP-element group 110: 	43 
    -- CP-element group 110: 	47 
    -- CP-element group 110: 	41 
    -- CP-element group 110: 	42 
    -- CP-element group 110:  members (33) 
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/word_access_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/word_access_complete/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/ptr_deref_1560_Update/word_access_complete/word_0/cr
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_update_start
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_complete/req
      -- CP-element group 110: 	 branch_block_stmt_1278/merge_stmt_1507__exit__
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563__entry__
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1511_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/addr_of_1557_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1550_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Update/req
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/array_obj_ref_1556_final_index_sum_regn_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/assign_stmt_1512_to_assign_stmt_1563/type_cast_1516_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1278/merge_stmt_1507_PhiReqMerge
      -- CP-element group 110: 	 branch_block_stmt_1278/merge_stmt_1507_PhiAck/$entry
      -- CP-element group 110: 	 branch_block_stmt_1278/merge_stmt_1507_PhiAck/$exit
      -- CP-element group 110: 	 branch_block_stmt_1278/merge_stmt_1507_PhiAck/dummy
      -- 
    rr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => type_cast_1511_inst_req_0); -- 
    cr_4047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => ptr_deref_1560_store_0_req_1); -- 
    cr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => type_cast_1550_inst_req_1); -- 
    cr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => type_cast_1511_inst_req_1); -- 
    req_3997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => addr_of_1557_final_reg_req_1); -- 
    cr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => type_cast_1516_inst_req_1); -- 
    req_3982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => array_obj_ref_1556_index_offset_req_1); -- 
    rr_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(110), ack => type_cast_1516_inst_req_0); -- 
    zeropad3D_B_CP_3564_elements(110) <= OrReduce(zeropad3D_B_CP_3564_elements(36) & zeropad3D_B_CP_3564_elements(40));
    -- CP-element group 111:  merge  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	54 
    -- CP-element group 111: 	74 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	75 
    -- CP-element group 111: 	76 
    -- CP-element group 111:  members (13) 
      -- CP-element group 111: 	 branch_block_stmt_1278/merge_stmt_1672__exit__
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690__entry__
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/$entry
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1278/assign_stmt_1677_to_assign_stmt_1690/type_cast_1676_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_1278/merge_stmt_1672_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_1278/merge_stmt_1672_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_1278/merge_stmt_1672_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_1278/merge_stmt_1672_PhiAck/dummy
      -- 
    rr_4296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(111), ack => type_cast_1676_inst_req_0); -- 
    cr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(111), ack => type_cast_1676_inst_req_1); -- 
    zeropad3D_B_CP_3564_elements(111) <= OrReduce(zeropad3D_B_CP_3564_elements(54) & zeropad3D_B_CP_3564_elements(74));
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Sample/ra
      -- 
    ra_4616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1766_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/Update/ca
      -- 
    ca_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1766_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	119 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/$exit
      -- CP-element group 114: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/$exit
      -- CP-element group 114: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1766/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_req
      -- 
    phi_stmt_1761_req_4622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1761_req_4622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(114), ack => phi_stmt_1761_req_1); -- 
    zeropad3D_B_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(112) & zeropad3D_B_CP_3564_elements(113);
      gj_zeropad3D_B_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	86 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Sample/ra
      -- 
    ra_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/Update/ca
      -- 
    ca_4644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/$exit
      -- CP-element group 117: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/$exit
      -- CP-element group 117: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1772/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_req
      -- 
    phi_stmt_1767_req_4645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1767_req_4645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(117), ack => phi_stmt_1767_req_1); -- 
    zeropad3D_B_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(115) & zeropad3D_B_CP_3564_elements(116);
      gj_zeropad3D_B_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  output  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	86 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1754/$exit
      -- CP-element group 118: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1760_konst_delay_trans
      -- CP-element group 118: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_req
      -- 
    phi_stmt_1754_req_4653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1754_req_4653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(118), ack => phi_stmt_1754_req_1); -- 
    -- Element group zeropad3D_B_CP_3564_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_3564_elements(86), ack => zeropad3D_B_CP_3564_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  join  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	114 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	130 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1278/ifx_xelse151_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(114) & zeropad3D_B_CP_3564_elements(117) & zeropad3D_B_CP_3564_elements(118);
      gj_zeropad3D_B_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Sample/ra
      -- 
    ra_4673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/Update/ca
      -- 
    ca_4678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	129 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/$exit
      -- CP-element group 122: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/$exit
      -- CP-element group 122: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_sources/type_cast_1764/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1761/phi_stmt_1761_req
      -- 
    phi_stmt_1761_req_4679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1761_req_4679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(122), ack => phi_stmt_1761_req_0); -- 
    zeropad3D_B_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(120) & zeropad3D_B_CP_3564_elements(121);
      gj_zeropad3D_B_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Sample/ra
      -- 
    ra_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1770_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/Update/ca
      -- 
    ca_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1770_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/$exit
      -- CP-element group 125: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/$exit
      -- CP-element group 125: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_sources/type_cast_1770/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1767/phi_stmt_1767_req
      -- 
    phi_stmt_1767_req_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1767_req_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(125), ack => phi_stmt_1767_req_0); -- 
    zeropad3D_B_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(123) & zeropad3D_B_CP_3564_elements(124);
      gj_zeropad3D_B_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Sample/ra
      -- 
    ra_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1757_inst_ack_0, ack => zeropad3D_B_CP_3564_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	77 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/Update/ca
      -- 
    ca_4724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1757_inst_ack_1, ack => zeropad3D_B_CP_3564_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/$exit
      -- CP-element group 128: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/$exit
      -- CP-element group 128: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/type_cast_1757/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1754/phi_stmt_1754_req
      -- 
    phi_stmt_1754_req_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1754_req_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3564_elements(128), ack => phi_stmt_1754_req_0); -- 
    zeropad3D_B_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(126) & zeropad3D_B_CP_3564_elements(127);
      gj_zeropad3D_B_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1278/ifx_xthen146_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(122) & zeropad3D_B_CP_3564_elements(125) & zeropad3D_B_CP_3564_elements(128);
      gj_zeropad3D_B_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1278/merge_stmt_1753_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1278/merge_stmt_1753_PhiAck/$entry
      -- 
    zeropad3D_B_CP_3564_elements(130) <= OrReduce(zeropad3D_B_CP_3564_elements(119) & zeropad3D_B_CP_3564_elements(129));
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1278/merge_stmt_1753_PhiAck/phi_stmt_1754_ack
      -- 
    phi_stmt_1754_ack_4730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1754_ack_0, ack => zeropad3D_B_CP_3564_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1278/merge_stmt_1753_PhiAck/phi_stmt_1761_ack
      -- 
    phi_stmt_1761_ack_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1761_ack_0, ack => zeropad3D_B_CP_3564_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1278/merge_stmt_1753_PhiAck/phi_stmt_1767_ack
      -- 
    phi_stmt_1767_ack_4732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1767_ack_0, ack => zeropad3D_B_CP_3564_elements(133)); -- 
    -- CP-element group 134:  join  transition  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	1 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1278/merge_stmt_1753_PhiAck/$exit
      -- 
    zeropad3D_B_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3564_elements(131) & zeropad3D_B_CP_3564_elements(132) & zeropad3D_B_CP_3564_elements(133);
      gj_zeropad3D_B_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3564_elements(134), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1352_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1408_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1544_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1627_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1652_wire : std_logic_vector(31 downto 0);
    signal R_idxprom131_1638_resized : std_logic_vector(13 downto 0);
    signal R_idxprom131_1638_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom136_1663_resized : std_logic_vector(13 downto 0);
    signal R_idxprom136_1663_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1555_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1555_scaled : std_logic_vector(13 downto 0);
    signal add103_1595 : std_logic_vector(31 downto 0);
    signal add112_1600 : std_logic_vector(31 downto 0);
    signal add122_1615 : std_logic_vector(31 downto 0);
    signal add128_1620 : std_logic_vector(31 downto 0);
    signal add141_1683 : std_logic_vector(31 downto 0);
    signal add149_1703 : std_logic_vector(15 downto 0);
    signal add159_1365 : std_logic_vector(31 downto 0);
    signal add175_1380 : std_logic_vector(31 downto 0);
    signal add74_1390 : std_logic_vector(31 downto 0);
    signal add85_1532 : std_logic_vector(31 downto 0);
    signal add91_1537 : std_logic_vector(31 downto 0);
    signal add_1385 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1556_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1556_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1556_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1556_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1556_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1556_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1639_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1639_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1639_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1639_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1639_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1639_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1664_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1664_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1664_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1664_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1664_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1664_root_address : std_logic_vector(13 downto 0);
    signal arrayidx132_1641 : std_logic_vector(31 downto 0);
    signal arrayidx137_1666 : std_logic_vector(31 downto 0);
    signal arrayidx_1558 : std_logic_vector(31 downto 0);
    signal call1_1284 : std_logic_vector(7 downto 0);
    signal call2_1287 : std_logic_vector(7 downto 0);
    signal call3_1290 : std_logic_vector(7 downto 0);
    signal call4_1293 : std_logic_vector(7 downto 0);
    signal call5_1296 : std_logic_vector(7 downto 0);
    signal call6_1299 : std_logic_vector(7 downto 0);
    signal call_1281 : std_logic_vector(7 downto 0);
    signal cmp144_1690 : std_logic_vector(0 downto 0);
    signal cmp160_1721 : std_logic_vector(0 downto 0);
    signal cmp176_1746 : std_logic_vector(0 downto 0);
    signal cmp58_1458 : std_logic_vector(0 downto 0);
    signal cmp65_1482 : std_logic_vector(0 downto 0);
    signal cmp65x_xnot_1488 : std_logic_vector(0 downto 0);
    signal cmp75_1495 : std_logic_vector(0 downto 0);
    signal cmp_1445 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_1451 : std_logic_vector(0 downto 0);
    signal conv105_1410 : std_logic_vector(31 downto 0);
    signal conv140_1677 : std_logic_vector(31 downto 0);
    signal conv154_1716 : std_logic_vector(31 downto 0);
    signal conv168_1741 : std_logic_vector(31 downto 0);
    signal conv170_1369 : std_logic_vector(31 downto 0);
    signal conv32_1314 : std_logic_vector(31 downto 0);
    signal conv34_1318 : std_logic_vector(31 downto 0);
    signal conv38_1322 : std_logic_vector(31 downto 0);
    signal conv40_1326 : std_logic_vector(31 downto 0);
    signal conv47_1438 : std_logic_vector(31 downto 0);
    signal conv49_1335 : std_logic_vector(31 downto 0);
    signal conv62_1475 : std_logic_vector(31 downto 0);
    signal conv79_1512 : std_logic_vector(31 downto 0);
    signal conv81_1339 : std_logic_vector(31 downto 0);
    signal conv83_1517 : std_logic_vector(31 downto 0);
    signal conv87_1354 : std_logic_vector(31 downto 0);
    signal conv95_1570 : std_logic_vector(31 downto 0);
    signal conv_1304 : std_logic_vector(15 downto 0);
    signal div171_1375 : std_logic_vector(31 downto 0);
    signal div_1310 : std_logic_vector(15 downto 0);
    signal idxprom131_1634 : std_logic_vector(63 downto 0);
    signal idxprom136_1659 : std_logic_vector(63 downto 0);
    signal idxprom_1551 : std_logic_vector(63 downto 0);
    signal inc165_1725 : std_logic_vector(15 downto 0);
    signal inc165x_xix_x2_1730 : std_logic_vector(15 downto 0);
    signal inc_1711 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1761 : std_logic_vector(15 downto 0);
    signal ix_x2_1420 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1767 : std_logic_vector(15 downto 0);
    signal jx_x1_1427 : std_logic_vector(15 downto 0);
    signal jx_x2_1736 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1754 : std_logic_vector(15 downto 0);
    signal kx_x1_1413 : std_logic_vector(15 downto 0);
    signal mul102_1580 : std_logic_vector(31 downto 0);
    signal mul111_1590 : std_logic_vector(31 downto 0);
    signal mul121_1605 : std_logic_vector(31 downto 0);
    signal mul127_1610 : std_logic_vector(31 downto 0);
    signal mul41_1331 : std_logic_vector(31 downto 0);
    signal mul84_1522 : std_logic_vector(31 downto 0);
    signal mul90_1527 : std_logic_vector(31 downto 0);
    signal mul_1396 : std_logic_vector(31 downto 0);
    signal orx_xcond190_1500 : std_logic_vector(0 downto 0);
    signal orx_xcond_1463 : std_logic_vector(0 downto 0);
    signal ptr_deref_1560_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1560_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1560_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1560_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1560_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1560_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1644_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1644_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1644_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1644_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1644_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1668_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1668_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1668_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1668_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1668_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1668_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext189_1345 : std_logic_vector(31 downto 0);
    signal sext_1401 : std_logic_vector(31 downto 0);
    signal shl_1360 : std_logic_vector(31 downto 0);
    signal shr130_1629 : std_logic_vector(31 downto 0);
    signal shr135_1654 : std_logic_vector(31 downto 0);
    signal shr_1546 : std_logic_vector(31 downto 0);
    signal sub110_1585 : std_logic_vector(31 downto 0);
    signal sub_1575 : std_logic_vector(31 downto 0);
    signal tmp133_1645 : std_logic_vector(63 downto 0);
    signal type_cast_1308_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1343_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1348_wire : std_logic_vector(31 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1358_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1373_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1404_wire : std_logic_vector(31 downto 0);
    signal type_cast_1407_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1417_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1419_wire : std_logic_vector(15 downto 0);
    signal type_cast_1424_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1426_wire : std_logic_vector(15 downto 0);
    signal type_cast_1430_wire : std_logic_vector(15 downto 0);
    signal type_cast_1432_wire : std_logic_vector(15 downto 0);
    signal type_cast_1436_wire : std_logic_vector(31 downto 0);
    signal type_cast_1441_wire : std_logic_vector(31 downto 0);
    signal type_cast_1443_wire : std_logic_vector(31 downto 0);
    signal type_cast_1449_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1454_wire : std_logic_vector(31 downto 0);
    signal type_cast_1456_wire : std_logic_vector(31 downto 0);
    signal type_cast_1473_wire : std_logic_vector(31 downto 0);
    signal type_cast_1478_wire : std_logic_vector(31 downto 0);
    signal type_cast_1480_wire : std_logic_vector(31 downto 0);
    signal type_cast_1486_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1491_wire : std_logic_vector(31 downto 0);
    signal type_cast_1493_wire : std_logic_vector(31 downto 0);
    signal type_cast_1510_wire : std_logic_vector(31 downto 0);
    signal type_cast_1515_wire : std_logic_vector(31 downto 0);
    signal type_cast_1540_wire : std_logic_vector(31 downto 0);
    signal type_cast_1543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1549_wire : std_logic_vector(63 downto 0);
    signal type_cast_1562_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1568_wire : std_logic_vector(31 downto 0);
    signal type_cast_1623_wire : std_logic_vector(31 downto 0);
    signal type_cast_1626_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1632_wire : std_logic_vector(63 downto 0);
    signal type_cast_1648_wire : std_logic_vector(31 downto 0);
    signal type_cast_1651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1657_wire : std_logic_vector(63 downto 0);
    signal type_cast_1675_wire : std_logic_vector(31 downto 0);
    signal type_cast_1681_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1686_wire : std_logic_vector(31 downto 0);
    signal type_cast_1688_wire : std_logic_vector(31 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1709_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1714_wire : std_logic_vector(31 downto 0);
    signal type_cast_1739_wire : std_logic_vector(31 downto 0);
    signal type_cast_1757_wire : std_logic_vector(15 downto 0);
    signal type_cast_1760_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1764_wire : std_logic_vector(15 downto 0);
    signal type_cast_1766_wire : std_logic_vector(15 downto 0);
    signal type_cast_1770_wire : std_logic_vector(15 downto 0);
    signal type_cast_1772_wire : std_logic_vector(15 downto 0);
    signal type_cast_1779_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1556_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1556_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1556_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1556_resized_base_address <= "00000000000000";
    array_obj_ref_1639_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1639_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1639_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1639_resized_base_address <= "00000000000000";
    array_obj_ref_1664_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1664_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1664_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1664_resized_base_address <= "00000000000000";
    ptr_deref_1560_word_offset_0 <= "00000000000000";
    ptr_deref_1644_word_offset_0 <= "00000000000000";
    ptr_deref_1668_word_offset_0 <= "00000000000000";
    type_cast_1308_wire_constant <= "0000000000000001";
    type_cast_1343_wire_constant <= "00000000000000000000000000010000";
    type_cast_1351_wire_constant <= "00000000000000000000000000010000";
    type_cast_1358_wire_constant <= "00000000000000000000000000000001";
    type_cast_1373_wire_constant <= "00000000000000000000000000000010";
    type_cast_1394_wire_constant <= "00000000000000000000000000010000";
    type_cast_1407_wire_constant <= "00000000000000000000000000010000";
    type_cast_1417_wire_constant <= "0000000000000000";
    type_cast_1424_wire_constant <= "0000000000000000";
    type_cast_1449_wire_constant <= "1";
    type_cast_1486_wire_constant <= "1";
    type_cast_1543_wire_constant <= "00000000000000000000000000000010";
    type_cast_1562_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1626_wire_constant <= "00000000000000000000000000000010";
    type_cast_1651_wire_constant <= "00000000000000000000000000000010";
    type_cast_1681_wire_constant <= "00000000000000000000000000000100";
    type_cast_1701_wire_constant <= "0000000000000100";
    type_cast_1709_wire_constant <= "0000000000000001";
    type_cast_1760_wire_constant <= "0000000000000000";
    type_cast_1779_wire_constant <= "00000001";
    phi_stmt_1413: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1417_wire_constant & type_cast_1419_wire;
      req <= phi_stmt_1413_req_0 & phi_stmt_1413_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1413",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1413_ack_0,
          idata => idata,
          odata => kx_x1_1413,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1413
    phi_stmt_1420: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1424_wire_constant & type_cast_1426_wire;
      req <= phi_stmt_1420_req_0 & phi_stmt_1420_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1420",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1420_ack_0,
          idata => idata,
          odata => ix_x2_1420,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1420
    phi_stmt_1427: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1430_wire & type_cast_1432_wire;
      req <= phi_stmt_1427_req_0 & phi_stmt_1427_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1427",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1427_ack_0,
          idata => idata,
          odata => jx_x1_1427,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1427
    phi_stmt_1754: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1757_wire & type_cast_1760_wire_constant;
      req <= phi_stmt_1754_req_0 & phi_stmt_1754_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1754",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1754_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1754,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1754
    phi_stmt_1761: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1764_wire & type_cast_1766_wire;
      req <= phi_stmt_1761_req_0 & phi_stmt_1761_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1761",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1761_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1761,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1761
    phi_stmt_1767: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1770_wire & type_cast_1772_wire;
      req <= phi_stmt_1767_req_0 & phi_stmt_1767_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1767",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1767_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1767,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1767
    -- flow-through select operator MUX_1735_inst
    jx_x2_1736 <= div_1310 when (cmp160_1721(0) /=  '0') else inc_1711;
    addr_of_1557_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1557_final_reg_req_0;
      addr_of_1557_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1557_final_reg_req_1;
      addr_of_1557_final_reg_ack_1<= rack(0);
      addr_of_1557_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1557_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1556_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1640_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1640_final_reg_req_0;
      addr_of_1640_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1640_final_reg_req_1;
      addr_of_1640_final_reg_ack_1<= rack(0);
      addr_of_1640_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1640_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1639_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx132_1641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1665_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1665_final_reg_req_0;
      addr_of_1665_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1665_final_reg_req_1;
      addr_of_1665_final_reg_ack_1<= rack(0);
      addr_of_1665_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1665_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1664_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx137_1666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1303_inst_req_0;
      type_cast_1303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1303_inst_req_1;
      type_cast_1303_inst_ack_1<= rack(0);
      type_cast_1303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1313_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1313_inst_req_0;
      type_cast_1313_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1313_inst_req_1;
      type_cast_1313_inst_ack_1<= rack(0);
      type_cast_1313_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1313_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1314,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1317_inst_req_0;
      type_cast_1317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1317_inst_req_1;
      type_cast_1317_inst_ack_1<= rack(0);
      type_cast_1317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_1318,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1321_inst_req_0;
      type_cast_1321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1321_inst_req_1;
      type_cast_1321_inst_ack_1<= rack(0);
      type_cast_1321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_1322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1325_inst_req_0;
      type_cast_1325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1325_inst_req_1;
      type_cast_1325_inst_ack_1<= rack(0);
      type_cast_1325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_1293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_1326,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1334_inst_req_0;
      type_cast_1334_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1334_inst_req_1;
      type_cast_1334_inst_ack_1<= rack(0);
      type_cast_1334_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1334_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1338_inst_req_0;
      type_cast_1338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1338_inst_req_1;
      type_cast_1338_inst_ack_1<= rack(0);
      type_cast_1338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1348_inst
    process(sext189_1345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext189_1345(31 downto 0);
      type_cast_1348_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1353_inst
    process(ASHR_i32_i32_1352_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1352_wire(31 downto 0);
      conv87_1354 <= tmp_var; -- 
    end process;
    type_cast_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1368_inst_req_0;
      type_cast_1368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1368_inst_req_1;
      type_cast_1368_inst_ack_1<= rack(0);
      type_cast_1368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1404_inst
    process(sext_1401) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1401(31 downto 0);
      type_cast_1404_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1409_inst
    process(ASHR_i32_i32_1408_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1408_wire(31 downto 0);
      conv105_1410 <= tmp_var; -- 
    end process;
    type_cast_1419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1419_inst_req_0;
      type_cast_1419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1419_inst_req_1;
      type_cast_1419_inst_ack_1<= rack(0);
      type_cast_1419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1419_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1426_inst_req_0;
      type_cast_1426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1426_inst_req_1;
      type_cast_1426_inst_ack_1<= rack(0);
      type_cast_1426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1426_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1430_inst_req_0;
      type_cast_1430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1430_inst_req_1;
      type_cast_1430_inst_ack_1<= rack(0);
      type_cast_1430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1430_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1432_inst_req_0;
      type_cast_1432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1432_inst_req_1;
      type_cast_1432_inst_ack_1<= rack(0);
      type_cast_1432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1437_inst_req_0;
      type_cast_1437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1437_inst_req_1;
      type_cast_1437_inst_ack_1<= rack(0);
      type_cast_1437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1436_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1441_inst
    process(conv47_1438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_1438(31 downto 0);
      type_cast_1441_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1443_inst
    process(conv49_1335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_1335(31 downto 0);
      type_cast_1443_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1454_inst
    process(conv47_1438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_1438(31 downto 0);
      type_cast_1454_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1456_inst
    process(add_1385) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_1385(31 downto 0);
      type_cast_1456_wire <= tmp_var; -- 
    end process;
    type_cast_1474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1474_inst_req_0;
      type_cast_1474_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1474_inst_req_1;
      type_cast_1474_inst_ack_1<= rack(0);
      type_cast_1474_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1474_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1473_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1478_inst
    process(conv62_1475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv62_1475(31 downto 0);
      type_cast_1478_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1480_inst
    process(conv49_1335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_1335(31 downto 0);
      type_cast_1480_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1491_inst
    process(conv62_1475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv62_1475(31 downto 0);
      type_cast_1491_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1493_inst
    process(add74_1390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add74_1390(31 downto 0);
      type_cast_1493_wire <= tmp_var; -- 
    end process;
    type_cast_1511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1511_inst_req_0;
      type_cast_1511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1511_inst_req_1;
      type_cast_1511_inst_ack_1<= rack(0);
      type_cast_1511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1510_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1516_inst_req_0;
      type_cast_1516_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1516_inst_req_1;
      type_cast_1516_inst_ack_1<= rack(0);
      type_cast_1516_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1516_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1515_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1517,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1540_inst
    process(add91_1537) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add91_1537(31 downto 0);
      type_cast_1540_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1545_inst
    process(ASHR_i32_i32_1544_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1544_wire(31 downto 0);
      shr_1546 <= tmp_var; -- 
    end process;
    type_cast_1550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1550_inst_req_0;
      type_cast_1550_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1550_inst_req_1;
      type_cast_1550_inst_ack_1<= rack(0);
      type_cast_1550_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1550_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1549_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1569_inst_req_0;
      type_cast_1569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1569_inst_req_1;
      type_cast_1569_inst_ack_1<= rack(0);
      type_cast_1569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1568_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_1570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1623_inst
    process(add112_1600) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add112_1600(31 downto 0);
      type_cast_1623_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1628_inst
    process(ASHR_i32_i32_1627_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1627_wire(31 downto 0);
      shr130_1629 <= tmp_var; -- 
    end process;
    type_cast_1633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1633_inst_req_0;
      type_cast_1633_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1633_inst_req_1;
      type_cast_1633_inst_ack_1<= rack(0);
      type_cast_1633_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1633_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1632_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom131_1634,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1648_inst
    process(add128_1620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add128_1620(31 downto 0);
      type_cast_1648_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1653_inst
    process(ASHR_i32_i32_1652_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1652_wire(31 downto 0);
      shr135_1654 <= tmp_var; -- 
    end process;
    type_cast_1658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1658_inst_req_0;
      type_cast_1658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1658_inst_req_1;
      type_cast_1658_inst_ack_1<= rack(0);
      type_cast_1658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1657_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom136_1659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1676_inst_req_0;
      type_cast_1676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1676_inst_req_1;
      type_cast_1676_inst_ack_1<= rack(0);
      type_cast_1676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1675_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_1677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1686_inst
    process(add141_1683) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add141_1683(31 downto 0);
      type_cast_1686_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1688_inst
    process(conv32_1314) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv32_1314(31 downto 0);
      type_cast_1688_wire <= tmp_var; -- 
    end process;
    type_cast_1715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1715_inst_req_0;
      type_cast_1715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1715_inst_req_1;
      type_cast_1715_inst_ack_1<= rack(0);
      type_cast_1715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1714_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_1716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1724_inst_req_0;
      type_cast_1724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1724_inst_req_1;
      type_cast_1724_inst_ack_1<= rack(0);
      type_cast_1724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp160_1721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc165_1725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1740_inst_req_0;
      type_cast_1740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1740_inst_req_1;
      type_cast_1740_inst_ack_1<= rack(0);
      type_cast_1740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1739_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv168_1741,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1757_inst_req_0;
      type_cast_1757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1757_inst_req_1;
      type_cast_1757_inst_ack_1<= rack(0);
      type_cast_1757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add149_1703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1757_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1764_inst_req_0;
      type_cast_1764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1764_inst_req_1;
      type_cast_1764_inst_ack_1<= rack(0);
      type_cast_1764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_1420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1764_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1766_inst_req_0;
      type_cast_1766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1766_inst_req_1;
      type_cast_1766_inst_ack_1<= rack(0);
      type_cast_1766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc165x_xix_x2_1730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1766_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1770_inst_req_0;
      type_cast_1770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1770_inst_req_1;
      type_cast_1770_inst_ack_1<= rack(0);
      type_cast_1770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_1427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1770_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1772_inst_req_0;
      type_cast_1772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1772_inst_req_1;
      type_cast_1772_inst_ack_1<= rack(0);
      type_cast_1772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1736,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1772_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1556_index_1_rename
    process(R_idxprom_1555_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1555_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1555_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1556_index_1_resize
    process(idxprom_1551) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1551;
      ov := iv(13 downto 0);
      R_idxprom_1555_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1556_root_address_inst
    process(array_obj_ref_1556_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1556_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1556_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1639_index_1_rename
    process(R_idxprom131_1638_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom131_1638_resized;
      ov(13 downto 0) := iv;
      R_idxprom131_1638_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1639_index_1_resize
    process(idxprom131_1634) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom131_1634;
      ov := iv(13 downto 0);
      R_idxprom131_1638_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1639_root_address_inst
    process(array_obj_ref_1639_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1639_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1639_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1664_index_1_rename
    process(R_idxprom136_1663_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom136_1663_resized;
      ov(13 downto 0) := iv;
      R_idxprom136_1663_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1664_index_1_resize
    process(idxprom136_1659) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom136_1659;
      ov := iv(13 downto 0);
      R_idxprom136_1663_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1664_root_address_inst
    process(array_obj_ref_1664_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1664_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1664_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1560_addr_0
    process(ptr_deref_1560_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1560_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1560_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1560_base_resize
    process(arrayidx_1558) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1558;
      ov := iv(13 downto 0);
      ptr_deref_1560_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1560_gather_scatter
    process(type_cast_1562_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1562_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1560_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1560_root_address_inst
    process(ptr_deref_1560_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1560_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1560_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1644_addr_0
    process(ptr_deref_1644_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1644_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1644_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1644_base_resize
    process(arrayidx132_1641) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx132_1641;
      ov := iv(13 downto 0);
      ptr_deref_1644_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1644_gather_scatter
    process(ptr_deref_1644_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1644_data_0;
      ov(63 downto 0) := iv;
      tmp133_1645 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1644_root_address_inst
    process(ptr_deref_1644_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1644_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1644_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1668_addr_0
    process(ptr_deref_1668_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1668_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1668_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1668_base_resize
    process(arrayidx137_1666) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx137_1666;
      ov := iv(13 downto 0);
      ptr_deref_1668_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1668_gather_scatter
    process(tmp133_1645) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp133_1645;
      ov(63 downto 0) := iv;
      ptr_deref_1668_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1668_root_address_inst
    process(ptr_deref_1668_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1668_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1668_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1464_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_1463;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1464_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1464_branch_req_0,
          ack0 => if_stmt_1464_branch_ack_0,
          ack1 => if_stmt_1464_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1501_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond190_1500;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1501_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1501_branch_req_0,
          ack0 => if_stmt_1501_branch_ack_0,
          ack1 => if_stmt_1501_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1691_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp144_1690;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1691_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1691_branch_req_0,
          ack0 => if_stmt_1691_branch_ack_0,
          ack1 => if_stmt_1691_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1747_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp176_1746;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1747_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1747_branch_req_0,
          ack0 => if_stmt_1747_branch_ack_0,
          ack1 => if_stmt_1747_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1702_inst
    process(kx_x1_1413) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_1413, type_cast_1701_wire_constant, tmp_var);
      add149_1703 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1710_inst
    process(jx_x1_1427) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_1427, type_cast_1709_wire_constant, tmp_var);
      inc_1711 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1729_inst
    process(inc165_1725, ix_x2_1420) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc165_1725, ix_x2_1420, tmp_var);
      inc165x_xix_x2_1730 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1364_inst
    process(shl_1360, conv34_1318) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1360, conv34_1318, tmp_var);
      add159_1365 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1379_inst
    process(shl_1360, div171_1375) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1360, div171_1375, tmp_var);
      add175_1380 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1384_inst
    process(conv49_1335, div171_1375) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv49_1335, div171_1375, tmp_var);
      add_1385 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1389_inst
    process(conv49_1335, conv34_1318) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv49_1335, conv34_1318, tmp_var);
      add74_1390 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1531_inst
    process(mul90_1527, conv79_1512) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul90_1527, conv79_1512, tmp_var);
      add85_1532 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1536_inst
    process(add85_1532, mul84_1522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add85_1532, mul84_1522, tmp_var);
      add91_1537 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1594_inst
    process(mul111_1590, conv95_1570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul111_1590, conv95_1570, tmp_var);
      add103_1595 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1599_inst
    process(add103_1595, mul102_1580) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add103_1595, mul102_1580, tmp_var);
      add112_1600 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1614_inst
    process(mul127_1610, conv95_1570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul127_1610, conv95_1570, tmp_var);
      add122_1615 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1619_inst
    process(add122_1615, mul121_1605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add122_1615, mul121_1605, tmp_var);
      add128_1620 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1682_inst
    process(conv140_1677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv140_1677, type_cast_1681_wire_constant, tmp_var);
      add141_1683 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1462_inst
    process(cmpx_xnot_1451, cmp58_1458) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_1451, cmp58_1458, tmp_var);
      orx_xcond_1463 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1499_inst
    process(cmp65x_xnot_1488, cmp75_1495) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp65x_xnot_1488, cmp75_1495, tmp_var);
      orx_xcond190_1500 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1352_inst
    process(type_cast_1348_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1348_wire, type_cast_1351_wire_constant, tmp_var);
      ASHR_i32_i32_1352_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1408_inst
    process(type_cast_1404_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1404_wire, type_cast_1407_wire_constant, tmp_var);
      ASHR_i32_i32_1408_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1544_inst
    process(type_cast_1540_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1540_wire, type_cast_1543_wire_constant, tmp_var);
      ASHR_i32_i32_1544_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1627_inst
    process(type_cast_1623_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1623_wire, type_cast_1626_wire_constant, tmp_var);
      ASHR_i32_i32_1627_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1652_inst
    process(type_cast_1648_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1648_wire, type_cast_1651_wire_constant, tmp_var);
      ASHR_i32_i32_1652_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1720_inst
    process(conv154_1716, add159_1365) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv154_1716, add159_1365, tmp_var);
      cmp160_1721 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1745_inst
    process(conv168_1741, add175_1380) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv168_1741, add175_1380, tmp_var);
      cmp176_1746 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1309_inst
    process(conv_1304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_1304, type_cast_1308_wire_constant, tmp_var);
      div_1310 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1374_inst
    process(conv170_1369) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv170_1369, type_cast_1373_wire_constant, tmp_var);
      div171_1375 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1330_inst
    process(conv38_1322, conv40_1326) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv38_1322, conv40_1326, tmp_var);
      mul41_1331 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1400_inst
    process(mul_1396, conv32_1314) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1396, conv32_1314, tmp_var);
      sext_1401 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1521_inst
    process(conv83_1517, conv81_1339) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv83_1517, conv81_1339, tmp_var);
      mul84_1522 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1526_inst
    process(conv47_1438, conv87_1354) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv47_1438, conv87_1354, tmp_var);
      mul90_1527 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1579_inst
    process(sub_1575, conv32_1314) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1575, conv32_1314, tmp_var);
      mul102_1580 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1589_inst
    process(sub110_1585, conv105_1410) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub110_1585, conv105_1410, tmp_var);
      mul111_1590 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1604_inst
    process(conv62_1475, conv81_1339) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv62_1475, conv81_1339, tmp_var);
      mul121_1605 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1609_inst
    process(conv47_1438, conv87_1354) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv47_1438, conv87_1354, tmp_var);
      mul127_1610 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1344_inst
    process(mul41_1331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul41_1331, type_cast_1343_wire_constant, tmp_var);
      sext189_1345 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1359_inst
    process(conv49_1335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1335, type_cast_1358_wire_constant, tmp_var);
      shl_1360 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1395_inst
    process(conv34_1318) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv34_1318, type_cast_1394_wire_constant, tmp_var);
      mul_1396 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1444_inst
    process(type_cast_1441_wire, type_cast_1443_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1441_wire, type_cast_1443_wire, tmp_var);
      cmp_1445 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1457_inst
    process(type_cast_1454_wire, type_cast_1456_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1454_wire, type_cast_1456_wire, tmp_var);
      cmp58_1458 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1481_inst
    process(type_cast_1478_wire, type_cast_1480_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1478_wire, type_cast_1480_wire, tmp_var);
      cmp65_1482 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1494_inst
    process(type_cast_1491_wire, type_cast_1493_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1491_wire, type_cast_1493_wire, tmp_var);
      cmp75_1495 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1689_inst
    process(type_cast_1686_wire, type_cast_1688_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1686_wire, type_cast_1688_wire, tmp_var);
      cmp144_1690 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1574_inst
    process(conv62_1475, conv49_1335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv62_1475, conv49_1335, tmp_var);
      sub_1575 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1584_inst
    process(conv47_1438, conv49_1335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv47_1438, conv49_1335, tmp_var);
      sub110_1585 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1450_inst
    process(cmp_1445) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_1445, type_cast_1449_wire_constant, tmp_var);
      cmpx_xnot_1451 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1487_inst
    process(cmp65_1482) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp65_1482, type_cast_1486_wire_constant, tmp_var);
      cmp65x_xnot_1488 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_1556_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1555_scaled;
      array_obj_ref_1556_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1556_index_offset_req_0;
      array_obj_ref_1556_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1556_index_offset_req_1;
      array_obj_ref_1556_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_1639_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom131_1638_scaled;
      array_obj_ref_1639_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1639_index_offset_req_0;
      array_obj_ref_1639_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1639_index_offset_req_1;
      array_obj_ref_1639_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_1664_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom136_1663_scaled;
      array_obj_ref_1664_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1664_index_offset_req_0;
      array_obj_ref_1664_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1664_index_offset_req_1;
      array_obj_ref_1664_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- unary operator type_cast_1436_inst
    process(ix_x2_1420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_1420, tmp_var);
      type_cast_1436_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1473_inst
    process(jx_x1_1427) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1427, tmp_var);
      type_cast_1473_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1510_inst
    process(kx_x1_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1413, tmp_var);
      type_cast_1510_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1515_inst
    process(jx_x1_1427) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1427, tmp_var);
      type_cast_1515_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1549_inst
    process(shr_1546) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1546, tmp_var);
      type_cast_1549_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1568_inst
    process(kx_x1_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1413, tmp_var);
      type_cast_1568_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1632_inst
    process(shr130_1629) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr130_1629, tmp_var);
      type_cast_1632_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1657_inst
    process(shr135_1654) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr135_1654, tmp_var);
      type_cast_1657_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1675_inst
    process(kx_x1_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1413, tmp_var);
      type_cast_1675_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1714_inst
    process(inc_1711) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1711, tmp_var);
      type_cast_1714_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1739_inst
    process(inc165x_xix_x2_1730) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc165x_xix_x2_1730, tmp_var);
      type_cast_1739_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1644_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1644_load_0_req_0;
      ptr_deref_1644_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1644_load_0_req_1;
      ptr_deref_1644_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1644_word_address_0;
      ptr_deref_1644_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1560_store_0 ptr_deref_1668_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1560_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1668_store_0_req_0;
      ptr_deref_1560_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1668_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1560_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1668_store_0_req_1;
      ptr_deref_1560_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1668_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1560_word_address_0 & ptr_deref_1668_word_address_0;
      data_in <= ptr_deref_1560_data_0 & ptr_deref_1668_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_starting_1298_inst RPIPE_Block1_starting_1295_inst RPIPE_Block1_starting_1292_inst RPIPE_Block1_starting_1289_inst RPIPE_Block1_starting_1286_inst RPIPE_Block1_starting_1283_inst RPIPE_Block1_starting_1280_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block1_starting_1298_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_starting_1295_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_starting_1292_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_starting_1289_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_starting_1286_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_starting_1283_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_starting_1280_inst_req_0;
      RPIPE_Block1_starting_1298_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_starting_1295_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_starting_1292_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_starting_1289_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_starting_1286_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_starting_1283_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_starting_1280_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block1_starting_1298_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_starting_1295_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_starting_1292_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_starting_1289_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_starting_1286_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_starting_1283_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_starting_1280_inst_req_1;
      RPIPE_Block1_starting_1298_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_starting_1295_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_starting_1292_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_starting_1289_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_starting_1286_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_starting_1283_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_starting_1280_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call6_1299 <= data_out(55 downto 48);
      call5_1296 <= data_out(47 downto 40);
      call4_1293 <= data_out(39 downto 32);
      call3_1290 <= data_out(31 downto 24);
      call2_1287 <= data_out(23 downto 16);
      call1_1284 <= data_out(15 downto 8);
      call_1281 <= data_out(7 downto 0);
      Block1_starting_read_0_gI: SplitGuardInterface generic map(name => "Block1_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block1_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_starting_pipe_read_req(0),
          oack => Block1_starting_pipe_read_ack(0),
          odata => Block1_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_complete_1777_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_complete_1777_inst_req_0;
      WPIPE_Block1_complete_1777_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_complete_1777_inst_req_1;
      WPIPE_Block1_complete_1777_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1779_wire_constant;
      Block1_complete_write_0_gI: SplitGuardInterface generic map(name => "Block1_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_complete_pipe_write_req(0),
          oack => Block1_complete_pipe_write_ack(0),
          odata => Block1_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_B_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_C is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block2_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_C;
architecture zeropad3D_C_arch of zeropad3D_C is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_C_CP_4749_start: Boolean;
  signal zeropad3D_C_CP_4749_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_starting_1800_inst_req_1 : boolean;
  signal type_cast_1811_inst_req_1 : boolean;
  signal type_cast_1821_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1800_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1806_inst_req_0 : boolean;
  signal type_cast_1821_inst_ack_1 : boolean;
  signal type_cast_1842_inst_ack_1 : boolean;
  signal type_cast_1833_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1803_inst_req_1 : boolean;
  signal type_cast_1825_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1803_inst_req_0 : boolean;
  signal type_cast_1811_inst_ack_1 : boolean;
  signal type_cast_1846_inst_req_0 : boolean;
  signal type_cast_1825_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1800_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1806_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1806_inst_req_1 : boolean;
  signal type_cast_1821_inst_ack_0 : boolean;
  signal type_cast_1833_inst_ack_1 : boolean;
  signal type_cast_1811_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1803_inst_ack_1 : boolean;
  signal type_cast_1833_inst_ack_0 : boolean;
  signal type_cast_1829_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1806_inst_ack_1 : boolean;
  signal type_cast_1842_inst_req_1 : boolean;
  signal type_cast_1842_inst_req_0 : boolean;
  signal type_cast_1825_inst_req_0 : boolean;
  signal type_cast_1833_inst_req_0 : boolean;
  signal type_cast_1842_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1803_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1800_inst_req_0 : boolean;
  signal type_cast_1829_inst_req_0 : boolean;
  signal type_cast_1821_inst_req_0 : boolean;
  signal type_cast_1829_inst_ack_1 : boolean;
  signal phi_stmt_2269_req_1 : boolean;
  signal phi_stmt_2276_req_0 : boolean;
  signal type_cast_1882_inst_ack_1 : boolean;
  signal type_cast_1825_inst_ack_0 : boolean;
  signal type_cast_1882_inst_req_0 : boolean;
  signal type_cast_1811_inst_req_0 : boolean;
  signal type_cast_1846_inst_ack_0 : boolean;
  signal type_cast_1882_inst_ack_0 : boolean;
  signal type_cast_1882_inst_req_1 : boolean;
  signal type_cast_1846_inst_req_1 : boolean;
  signal type_cast_1846_inst_ack_1 : boolean;
  signal type_cast_1829_inst_ack_0 : boolean;
  signal type_cast_2281_inst_req_0 : boolean;
  signal type_cast_2281_inst_ack_0 : boolean;
  signal type_cast_2281_inst_req_1 : boolean;
  signal type_cast_2281_inst_ack_1 : boolean;
  signal phi_stmt_2276_req_1 : boolean;
  signal RPIPE_Block2_starting_1788_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1788_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1788_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1788_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1791_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1791_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1791_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1791_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1794_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1794_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1794_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1794_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1797_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1797_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1797_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1797_inst_ack_1 : boolean;
  signal type_cast_1951_inst_req_0 : boolean;
  signal type_cast_1951_inst_ack_0 : boolean;
  signal type_cast_1951_inst_req_1 : boolean;
  signal type_cast_1951_inst_ack_1 : boolean;
  signal if_stmt_1978_branch_req_0 : boolean;
  signal if_stmt_1978_branch_ack_1 : boolean;
  signal if_stmt_1978_branch_ack_0 : boolean;
  signal type_cast_1988_inst_req_0 : boolean;
  signal type_cast_1988_inst_ack_0 : boolean;
  signal type_cast_1988_inst_req_1 : boolean;
  signal type_cast_1988_inst_ack_1 : boolean;
  signal if_stmt_2015_branch_req_0 : boolean;
  signal if_stmt_2015_branch_ack_1 : boolean;
  signal if_stmt_2015_branch_ack_0 : boolean;
  signal type_cast_2025_inst_req_0 : boolean;
  signal type_cast_2025_inst_ack_0 : boolean;
  signal type_cast_2025_inst_req_1 : boolean;
  signal type_cast_2025_inst_ack_1 : boolean;
  signal type_cast_2030_inst_req_0 : boolean;
  signal type_cast_2030_inst_ack_0 : boolean;
  signal type_cast_2030_inst_req_1 : boolean;
  signal type_cast_2030_inst_ack_1 : boolean;
  signal type_cast_2064_inst_req_0 : boolean;
  signal type_cast_2064_inst_ack_0 : boolean;
  signal type_cast_2064_inst_req_1 : boolean;
  signal type_cast_2064_inst_ack_1 : boolean;
  signal array_obj_ref_2070_index_offset_req_0 : boolean;
  signal array_obj_ref_2070_index_offset_ack_0 : boolean;
  signal array_obj_ref_2070_index_offset_req_1 : boolean;
  signal array_obj_ref_2070_index_offset_ack_1 : boolean;
  signal addr_of_2071_final_reg_req_0 : boolean;
  signal addr_of_2071_final_reg_ack_0 : boolean;
  signal addr_of_2071_final_reg_req_1 : boolean;
  signal addr_of_2071_final_reg_ack_1 : boolean;
  signal ptr_deref_2074_store_0_req_0 : boolean;
  signal ptr_deref_2074_store_0_ack_0 : boolean;
  signal ptr_deref_2074_store_0_req_1 : boolean;
  signal ptr_deref_2074_store_0_ack_1 : boolean;
  signal type_cast_2083_inst_req_0 : boolean;
  signal type_cast_2083_inst_ack_0 : boolean;
  signal type_cast_2083_inst_req_1 : boolean;
  signal type_cast_2083_inst_ack_1 : boolean;
  signal type_cast_2147_inst_req_0 : boolean;
  signal type_cast_2147_inst_ack_0 : boolean;
  signal type_cast_2147_inst_req_1 : boolean;
  signal type_cast_2147_inst_ack_1 : boolean;
  signal type_cast_2272_inst_ack_0 : boolean;
  signal type_cast_2272_inst_req_0 : boolean;
  signal array_obj_ref_2153_index_offset_req_0 : boolean;
  signal phi_stmt_2282_ack_0 : boolean;
  signal array_obj_ref_2153_index_offset_ack_0 : boolean;
  signal array_obj_ref_2153_index_offset_req_1 : boolean;
  signal phi_stmt_2276_ack_0 : boolean;
  signal array_obj_ref_2153_index_offset_ack_1 : boolean;
  signal phi_stmt_2269_ack_0 : boolean;
  signal addr_of_2154_final_reg_req_0 : boolean;
  signal addr_of_2154_final_reg_ack_0 : boolean;
  signal phi_stmt_2282_req_0 : boolean;
  signal addr_of_2154_final_reg_req_1 : boolean;
  signal addr_of_2154_final_reg_ack_1 : boolean;
  signal type_cast_2285_inst_ack_1 : boolean;
  signal type_cast_2285_inst_req_1 : boolean;
  signal type_cast_2279_inst_ack_1 : boolean;
  signal type_cast_2279_inst_req_1 : boolean;
  signal ptr_deref_2158_load_0_req_0 : boolean;
  signal ptr_deref_2158_load_0_ack_0 : boolean;
  signal ptr_deref_2158_load_0_req_1 : boolean;
  signal ptr_deref_2158_load_0_ack_1 : boolean;
  signal type_cast_2172_inst_req_0 : boolean;
  signal type_cast_2172_inst_ack_0 : boolean;
  signal type_cast_2172_inst_req_1 : boolean;
  signal type_cast_2285_inst_ack_0 : boolean;
  signal type_cast_2172_inst_ack_1 : boolean;
  signal phi_stmt_2282_req_1 : boolean;
  signal phi_stmt_2269_req_0 : boolean;
  signal type_cast_2287_inst_ack_1 : boolean;
  signal type_cast_2287_inst_req_1 : boolean;
  signal array_obj_ref_2178_index_offset_req_0 : boolean;
  signal type_cast_2285_inst_req_0 : boolean;
  signal array_obj_ref_2178_index_offset_ack_0 : boolean;
  signal array_obj_ref_2178_index_offset_req_1 : boolean;
  signal array_obj_ref_2178_index_offset_ack_1 : boolean;
  signal addr_of_2179_final_reg_req_0 : boolean;
  signal addr_of_2179_final_reg_ack_0 : boolean;
  signal addr_of_2179_final_reg_req_1 : boolean;
  signal addr_of_2179_final_reg_ack_1 : boolean;
  signal type_cast_2287_inst_ack_0 : boolean;
  signal type_cast_2287_inst_req_0 : boolean;
  signal type_cast_2272_inst_ack_1 : boolean;
  signal type_cast_2279_inst_ack_0 : boolean;
  signal type_cast_2279_inst_req_0 : boolean;
  signal ptr_deref_2182_store_0_req_0 : boolean;
  signal ptr_deref_2182_store_0_ack_0 : boolean;
  signal type_cast_2272_inst_req_1 : boolean;
  signal ptr_deref_2182_store_0_req_1 : boolean;
  signal ptr_deref_2182_store_0_ack_1 : boolean;
  signal type_cast_2190_inst_req_0 : boolean;
  signal type_cast_2190_inst_ack_0 : boolean;
  signal type_cast_2190_inst_req_1 : boolean;
  signal type_cast_2190_inst_ack_1 : boolean;
  signal if_stmt_2205_branch_req_0 : boolean;
  signal if_stmt_2205_branch_ack_1 : boolean;
  signal if_stmt_2205_branch_ack_0 : boolean;
  signal type_cast_2229_inst_req_0 : boolean;
  signal type_cast_2229_inst_ack_0 : boolean;
  signal type_cast_2229_inst_req_1 : boolean;
  signal type_cast_2229_inst_ack_1 : boolean;
  signal type_cast_2238_inst_req_0 : boolean;
  signal type_cast_2238_inst_ack_0 : boolean;
  signal type_cast_2238_inst_req_1 : boolean;
  signal type_cast_2238_inst_ack_1 : boolean;
  signal type_cast_2255_inst_req_0 : boolean;
  signal type_cast_2255_inst_ack_0 : boolean;
  signal type_cast_2255_inst_req_1 : boolean;
  signal type_cast_2255_inst_ack_1 : boolean;
  signal if_stmt_2262_branch_req_0 : boolean;
  signal if_stmt_2262_branch_ack_1 : boolean;
  signal if_stmt_2262_branch_ack_0 : boolean;
  signal WPIPE_Block2_complete_2292_inst_req_0 : boolean;
  signal WPIPE_Block2_complete_2292_inst_ack_0 : boolean;
  signal WPIPE_Block2_complete_2292_inst_req_1 : boolean;
  signal WPIPE_Block2_complete_2292_inst_ack_1 : boolean;
  signal phi_stmt_1940_req_0 : boolean;
  signal type_cast_1937_inst_req_0 : boolean;
  signal type_cast_1937_inst_ack_0 : boolean;
  signal type_cast_1937_inst_req_1 : boolean;
  signal type_cast_1937_inst_ack_1 : boolean;
  signal phi_stmt_1934_req_0 : boolean;
  signal phi_stmt_1927_req_0 : boolean;
  signal type_cast_1946_inst_req_0 : boolean;
  signal type_cast_1946_inst_ack_0 : boolean;
  signal type_cast_1946_inst_req_1 : boolean;
  signal type_cast_1946_inst_ack_1 : boolean;
  signal phi_stmt_1940_req_1 : boolean;
  signal type_cast_1939_inst_req_0 : boolean;
  signal type_cast_1939_inst_ack_0 : boolean;
  signal type_cast_1939_inst_req_1 : boolean;
  signal type_cast_1939_inst_ack_1 : boolean;
  signal phi_stmt_1934_req_1 : boolean;
  signal type_cast_1933_inst_req_0 : boolean;
  signal type_cast_1933_inst_ack_0 : boolean;
  signal type_cast_1933_inst_req_1 : boolean;
  signal type_cast_1933_inst_ack_1 : boolean;
  signal phi_stmt_1927_req_1 : boolean;
  signal phi_stmt_1927_ack_0 : boolean;
  signal phi_stmt_1934_ack_0 : boolean;
  signal phi_stmt_1940_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_C_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_C_CP_4749_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_C_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_C_CP_4749_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_C_CP_4749_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_C_CP_4749_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_C_CP_4749: Block -- control-path 
    signal zeropad3D_C_CP_4749_elements: BooleanArray(134 downto 0);
    -- 
  begin -- 
    zeropad3D_C_CP_4749_elements(0) <= zeropad3D_C_CP_4749_start;
    zeropad3D_C_CP_4749_symbol <= zeropad3D_C_CP_4749_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1786/$entry
      -- CP-element group 0: 	 branch_block_stmt_1786/branch_block_stmt_1786__entry__
      -- CP-element group 0: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807__entry__
      -- CP-element group 0: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/$entry
      -- CP-element group 0: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Sample/rr
      -- 
    rr_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(0), ack => RPIPE_Block2_starting_1788_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	134 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	102 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_1786/merge_stmt_2268__exit__
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Update/cr
      -- 
    rr_5651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(1), ack => type_cast_1946_inst_req_0); -- 
    cr_5656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(1), ack => type_cast_1946_inst_req_1); -- 
    rr_5674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(1), ack => type_cast_1939_inst_req_0); -- 
    cr_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(1), ack => type_cast_1939_inst_req_1); -- 
    rr_5697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(1), ack => type_cast_1933_inst_req_0); -- 
    cr_5702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(1), ack => type_cast_1933_inst_req_1); -- 
    zeropad3D_C_CP_4749_elements(1) <= zeropad3D_C_CP_4749_elements(134);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Update/cr
      -- 
    ra_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1788_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(2)); -- 
    cr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(2), ack => RPIPE_Block2_starting_1788_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1788_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Sample/rr
      -- 
    ca_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1788_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(3)); -- 
    rr_4829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(3), ack => RPIPE_Block2_starting_1791_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Update/cr
      -- 
    ra_4830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1791_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(4)); -- 
    cr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(4), ack => RPIPE_Block2_starting_1791_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1791_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Sample/rr
      -- 
    ca_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1791_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(5)); -- 
    rr_4843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(5), ack => RPIPE_Block2_starting_1794_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Update/cr
      -- 
    ra_4844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1794_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(6)); -- 
    cr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(6), ack => RPIPE_Block2_starting_1794_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1794_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Sample/rr
      -- 
    ca_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1794_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(7)); -- 
    rr_4857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(7), ack => RPIPE_Block2_starting_1797_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Update/cr
      -- 
    ra_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1797_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(8)); -- 
    cr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(8), ack => RPIPE_Block2_starting_1797_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1797_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Sample/$entry
      -- 
    ca_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1797_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(9)); -- 
    rr_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(9), ack => RPIPE_Block2_starting_1800_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Sample/$exit
      -- 
    ra_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1800_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(10)); -- 
    cr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(10), ack => RPIPE_Block2_starting_1800_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1800_update_completed_
      -- 
    ca_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1800_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(11)); -- 
    rr_4885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(11), ack => RPIPE_Block2_starting_1803_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Sample/ra
      -- 
    ra_4886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1803_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(12)); -- 
    cr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(12), ack => RPIPE_Block2_starting_1803_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1803_update_completed_
      -- 
    ca_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1803_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(13)); -- 
    rr_4899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(13), ack => RPIPE_Block2_starting_1806_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_sample_completed_
      -- 
    ra_4900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1806_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(14)); -- 
    cr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(14), ack => RPIPE_Block2_starting_1806_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15:  members (55) 
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/RPIPE_Block2_starting_1806_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807__exit__
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924__entry__
      -- CP-element group 15: 	 branch_block_stmt_1786/assign_stmt_1789_to_assign_stmt_1807/$exit
      -- 
    ca_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1806_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(15)); -- 
    cr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1811_inst_req_1); -- 
    cr_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1821_inst_req_1); -- 
    cr_4977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1833_inst_req_1); -- 
    cr_4949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1825_inst_req_1); -- 
    rr_5000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1846_inst_req_0); -- 
    cr_4963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1829_inst_req_1); -- 
    cr_4991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1842_inst_req_1); -- 
    rr_4986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1842_inst_req_0); -- 
    rr_4944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1825_inst_req_0); -- 
    rr_4972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1833_inst_req_0); -- 
    rr_4958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1829_inst_req_0); -- 
    rr_4930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1821_inst_req_0); -- 
    rr_5014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1882_inst_req_0); -- 
    rr_4916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1811_inst_req_0); -- 
    cr_5019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1882_inst_req_1); -- 
    cr_5005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(15), ack => type_cast_1846_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Sample/$exit
      -- 
    ra_4917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1811_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1811_Update/$exit
      -- 
    ca_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1811_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Sample/ra
      -- 
    ra_4931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1821_update_completed_
      -- 
    ca_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Sample/ra
      -- 
    ra_4945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1825_update_completed_
      -- 
    ca_4950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Sample/ra
      -- 
    ra_4959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1829_Update/ca
      -- 
    ca_4964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Sample/ra
      -- 
    ra_4973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1833_update_completed_
      -- 
    ca_4978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_sample_completed_
      -- 
    ra_4987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1842_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1842_update_completed_
      -- 
    ca_4992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1842_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Sample/$exit
      -- 
    ra_5001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1846_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1846_Update/ca
      -- 
    ca_5006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1846_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Sample/ra
      -- 
    ra_5015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1882_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/type_cast_1882_update_completed_
      -- 
    ca_5020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1882_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	21 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	25 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: 	90 
    -- CP-element group 32: 	91 
    -- CP-element group 32: 	93 
    -- CP-element group 32:  members (16) 
      -- CP-element group 32: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924/$exit
      -- CP-element group 32: 	 branch_block_stmt_1786/assign_stmt_1812_to_assign_stmt_1924__exit__
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1940/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1927/$entry
      -- CP-element group 32: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/$entry
      -- 
    rr_5617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(32), ack => type_cast_1937_inst_req_0); -- 
    cr_5622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(32), ack => type_cast_1937_inst_req_1); -- 
    zeropad3D_C_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(31) & zeropad3D_C_CP_4749_elements(17) & zeropad3D_C_CP_4749_elements(19) & zeropad3D_C_CP_4749_elements(21) & zeropad3D_C_CP_4749_elements(23) & zeropad3D_C_CP_4749_elements(25) & zeropad3D_C_CP_4749_elements(27) & zeropad3D_C_CP_4749_elements(29);
      gj_zeropad3D_C_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	109 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Sample/ra
      -- 
    ra_5032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	109 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (13) 
      -- CP-element group 34: 	 branch_block_stmt_1786/R_orx_xcond_1979_place
      -- CP-element group 34: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/$exit
      -- CP-element group 34: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977__exit__
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978__entry__
      -- CP-element group 34: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978_eval_test/branch_req
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1786/if_stmt_1978_else_link/$entry
      -- 
    ca_5037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(34)); -- 
    branch_req_5045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(34), ack => if_stmt_1978_branch_req_0); -- 
    -- CP-element group 35:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (18) 
      -- CP-element group 35: 	 branch_block_stmt_1786/whilex_xbody_lorx_xlhsx_xfalse59
      -- CP-element group 35: 	 branch_block_stmt_1786/merge_stmt_1984__exit__
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014__entry__
      -- CP-element group 35: 	 branch_block_stmt_1786/if_stmt_1978_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_1786/if_stmt_1978_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/$entry
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1786/whilex_xbody_lorx_xlhsx_xfalse59_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_1786/whilex_xbody_lorx_xlhsx_xfalse59_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_1786/merge_stmt_1984_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_1786/merge_stmt_1984_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_1786/merge_stmt_1984_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_1786/merge_stmt_1984_PhiAck/dummy
      -- 
    if_choice_transition_5050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1978_branch_ack_1, ack => zeropad3D_C_CP_4749_elements(35)); -- 
    rr_5067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(35), ack => type_cast_1988_inst_req_0); -- 
    cr_5072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(35), ack => type_cast_1988_inst_req_1); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	110 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1786/whilex_xbody_ifx_xthen
      -- CP-element group 36: 	 branch_block_stmt_1786/if_stmt_1978_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_1786/if_stmt_1978_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_1786/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1786/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_5054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1978_branch_ack_0, ack => zeropad3D_C_CP_4749_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Sample/ra
      -- 
    ra_5068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1988_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (13) 
      -- CP-element group 38: 	 branch_block_stmt_1786/R_orx_xcond191_2016_place
      -- CP-element group 38: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014__exit__
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015__entry__
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015_else_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/$exit
      -- CP-element group 38: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1786/assign_stmt_1989_to_assign_stmt_2014/type_cast_1988_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015_eval_test/branch_req
      -- CP-element group 38: 	 branch_block_stmt_1786/if_stmt_2015_if_link/$entry
      -- 
    ca_5073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1988_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(38)); -- 
    branch_req_5081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(38), ack => if_stmt_2015_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_1786/lorx_xlhsx_xfalse59_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_1786/merge_stmt_2079__exit__
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184__entry__
      -- CP-element group 39: 	 branch_block_stmt_1786/if_stmt_2015_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_1786/if_stmt_2015_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1786/lorx_xlhsx_xfalse59_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/lorx_xlhsx_xfalse59_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_1786/merge_stmt_2079_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_1786/merge_stmt_2079_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_1786/merge_stmt_2079_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_1786/merge_stmt_2079_PhiAck/dummy
      -- 
    if_choice_transition_5086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2015_branch_ack_1, ack => zeropad3D_C_CP_4749_elements(39)); -- 
    rr_5244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => type_cast_2083_inst_req_0); -- 
    cr_5249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => type_cast_2083_inst_req_1); -- 
    cr_5263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => type_cast_2147_inst_req_1); -- 
    req_5294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => array_obj_ref_2153_index_offset_req_1); -- 
    req_5309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => addr_of_2154_final_reg_req_1); -- 
    cr_5354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => ptr_deref_2158_load_0_req_1); -- 
    cr_5373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => type_cast_2172_inst_req_1); -- 
    req_5404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => array_obj_ref_2178_index_offset_req_1); -- 
    req_5419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => addr_of_2179_final_reg_req_1); -- 
    cr_5469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(39), ack => ptr_deref_2182_store_0_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	110 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1786/if_stmt_2015_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_1786/if_stmt_2015_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_1786/lorx_xlhsx_xfalse59_ifx_xthen
      -- CP-element group 40: 	 branch_block_stmt_1786/lorx_xlhsx_xfalse59_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_1786/lorx_xlhsx_xfalse59_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2015_branch_ack_0, ack => zeropad3D_C_CP_4749_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	110 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Sample/ra
      -- 
    ra_5104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	110 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Update/ca
      -- 
    ca_5109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	110 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Sample/ra
      -- 
    ra_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Update/ca
      -- 
    ca_5123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Sample/rr
      -- 
    rr_5131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(45), ack => type_cast_2064_inst_req_0); -- 
    zeropad3D_C_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(44) & zeropad3D_C_CP_4749_elements(42);
      gj_zeropad3D_C_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Sample/ra
      -- 
    ra_5132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2064_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	110 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_computed_1
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Sample/req
      -- 
    ca_5137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2064_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(47)); -- 
    req_5162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(47), ack => array_obj_ref_2070_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Sample/ack
      -- 
    ack_5163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2070_index_offset_ack_0, ack => zeropad3D_C_CP_4749_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	110 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_request/req
      -- 
    ack_5168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2070_index_offset_ack_1, ack => zeropad3D_C_CP_4749_elements(49)); -- 
    req_5177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(49), ack => addr_of_2071_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_request/$exit
      -- CP-element group 50: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_request/ack
      -- 
    ack_5178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2071_final_reg_ack_0, ack => zeropad3D_C_CP_4749_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	110 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_word_addrgen/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/ptr_deref_2074_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/ptr_deref_2074_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/ptr_deref_2074_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/ptr_deref_2074_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/word_access_start/word_0/rr
      -- 
    ack_5183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2071_final_reg_ack_1, ack => zeropad3D_C_CP_4749_elements(51)); -- 
    rr_5221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(51), ack => ptr_deref_2074_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Sample/word_access_start/word_0/ra
      -- 
    ra_5222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2074_store_0_ack_0, ack => zeropad3D_C_CP_4749_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	110 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/word_access_complete/word_0/ca
      -- 
    ca_5233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2074_store_0_ack_1, ack => zeropad3D_C_CP_4749_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: 	48 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	111 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1786/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077__exit__
      -- CP-element group 54: 	 branch_block_stmt_1786/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/$exit
      -- CP-element group 54: 	 branch_block_stmt_1786/ifx_xthen_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_C_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(53) & zeropad3D_C_CP_4749_elements(48);
      gj_zeropad3D_C_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Sample/ra
      -- 
    ra_5245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2083_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2083_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Sample/rr
      -- 
    ca_5250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2083_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(56)); -- 
    rr_5258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(56), ack => type_cast_2147_inst_req_0); -- 
    rr_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(56), ack => type_cast_2172_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Sample/ra
      -- 
    ra_5259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2147_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Sample/req
      -- 
    ca_5264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(58)); -- 
    req_5289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(58), ack => array_obj_ref_2153_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Sample/ack
      -- 
    ack_5290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2153_index_offset_ack_0, ack => zeropad3D_C_CP_4749_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2153_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_request/req
      -- 
    ack_5295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2153_index_offset_ack_1, ack => zeropad3D_C_CP_4749_elements(60)); -- 
    req_5304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(60), ack => addr_of_2154_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_request/ack
      -- 
    ack_5305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2154_final_reg_ack_0, ack => zeropad3D_C_CP_4749_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2154_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/word_access_start/word_0/rr
      -- 
    ack_5310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2154_final_reg_ack_1, ack => zeropad3D_C_CP_4749_elements(62)); -- 
    rr_5343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(62), ack => ptr_deref_2158_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Sample/word_access_start/word_0/ra
      -- 
    ra_5344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2158_load_0_ack_0, ack => zeropad3D_C_CP_4749_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/ptr_deref_2158_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/ptr_deref_2158_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/ptr_deref_2158_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2158_Update/ptr_deref_2158_Merge/merge_ack
      -- 
    ca_5355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2158_load_0_ack_1, ack => zeropad3D_C_CP_4749_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Sample/ra
      -- 
    ra_5369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2172_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/type_cast_2172_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_computed_1
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Sample/req
      -- 
    ca_5374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2172_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(66)); -- 
    req_5399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(66), ack => array_obj_ref_2178_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Sample/ack
      -- 
    ack_5400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2178_index_offset_ack_0, ack => zeropad3D_C_CP_4749_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/array_obj_ref_2178_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_request/req
      -- 
    ack_5405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2178_index_offset_ack_1, ack => zeropad3D_C_CP_4749_elements(68)); -- 
    req_5414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(68), ack => addr_of_2179_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_request/ack
      -- 
    ack_5415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2179_final_reg_ack_0, ack => zeropad3D_C_CP_4749_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/addr_of_2179_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_word_addrgen/root_register_ack
      -- 
    ack_5420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2179_final_reg_ack_1, ack => zeropad3D_C_CP_4749_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/ptr_deref_2182_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/ptr_deref_2182_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/ptr_deref_2182_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/ptr_deref_2182_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/word_access_start/word_0/rr
      -- 
    rr_5458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(71), ack => ptr_deref_2182_store_0_req_0); -- 
    zeropad3D_C_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(64) & zeropad3D_C_CP_4749_elements(70);
      gj_zeropad3D_C_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Sample/word_access_start/word_0/ra
      -- 
    ra_5459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2182_store_0_ack_0, ack => zeropad3D_C_CP_4749_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/ptr_deref_2182_Update/word_access_complete/word_0/ca
      -- 
    ca_5470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2182_store_0_ack_1, ack => zeropad3D_C_CP_4749_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	111 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184__exit__
      -- CP-element group 74: 	 branch_block_stmt_1786/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_1786/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_1786/assign_stmt_2084_to_assign_stmt_2184/$exit
      -- CP-element group 74: 	 branch_block_stmt_1786/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(59) & zeropad3D_C_CP_4749_elements(67) & zeropad3D_C_CP_4749_elements(73);
      gj_zeropad3D_C_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	111 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Sample/ra
      -- 
    ra_5482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2190_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	111 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204__exit__
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205__entry__
      -- CP-element group 76: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/$exit
      -- CP-element group 76: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_1786/R_cmp144_2206_place
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1786/if_stmt_2205_else_link/$entry
      -- 
    ca_5487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2190_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(76)); -- 
    branch_req_5495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(76), ack => if_stmt_2205_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	127 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/merge_stmt_2211_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xend_ifx_xthen146_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/merge_stmt_2211__exit__
      -- CP-element group 77: 	 branch_block_stmt_1786/assign_stmt_2217__entry__
      -- CP-element group 77: 	 branch_block_stmt_1786/assign_stmt_2217__exit__
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/merge_stmt_2211_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/merge_stmt_2211_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/merge_stmt_2211_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xend_ifx_xthen146_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_1786/if_stmt_2205_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_1786/if_stmt_2205_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_1786/ifx_xend_ifx_xthen146
      -- CP-element group 77: 	 branch_block_stmt_1786/assign_stmt_2217/$entry
      -- CP-element group 77: 	 branch_block_stmt_1786/assign_stmt_2217/$exit
      -- 
    if_choice_transition_5500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2205_branch_ack_1, ack => zeropad3D_C_CP_4749_elements(77)); -- 
    rr_5880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(77), ack => type_cast_2281_inst_req_0); -- 
    cr_5885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(77), ack => type_cast_2281_inst_req_1); -- 
    rr_5857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(77), ack => type_cast_2272_inst_req_0); -- 
    cr_5908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(77), ack => type_cast_2285_inst_req_1); -- 
    rr_5903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(77), ack => type_cast_2285_inst_req_0); -- 
    cr_5862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(77), ack => type_cast_2272_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (24) 
      -- CP-element group 78: 	 branch_block_stmt_1786/merge_stmt_2219_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1786/merge_stmt_2219_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1786/merge_stmt_2219_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1786/merge_stmt_2219__exit__
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261__entry__
      -- CP-element group 78: 	 branch_block_stmt_1786/merge_stmt_2219_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/ifx_xend_ifx_xelse151_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1786/ifx_xend_ifx_xelse151_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/if_stmt_2205_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_1786/if_stmt_2205_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_1786/ifx_xend_ifx_xelse151
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Update/cr
      -- 
    else_choice_transition_5504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2205_branch_ack_0, ack => zeropad3D_C_CP_4749_elements(78)); -- 
    rr_5520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(78), ack => type_cast_2229_inst_req_0); -- 
    cr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(78), ack => type_cast_2229_inst_req_1); -- 
    cr_5539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(78), ack => type_cast_2238_inst_req_1); -- 
    cr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(78), ack => type_cast_2255_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Sample/ra
      -- 
    ra_5521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2229_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2229_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Sample/rr
      -- 
    ca_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2229_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(80)); -- 
    rr_5534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(80), ack => type_cast_2238_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Sample/ra
      -- 
    ra_5535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2238_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Sample/rr
      -- 
    ca_5540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(82)); -- 
    rr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(82), ack => type_cast_2255_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Sample/ra
      -- 
    ra_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2255_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(83)); -- 
    -- CP-element group 84:  branch  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (13) 
      -- CP-element group 84: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261__exit__
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262__entry__
      -- CP-element group 84: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/$exit
      -- CP-element group 84: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1786/assign_stmt_2225_to_assign_stmt_2261/type_cast_2255_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_1786/R_cmp177_2263_place
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1786/if_stmt_2262_else_link/$entry
      -- 
    ca_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2255_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(84)); -- 
    branch_req_5562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(84), ack => if_stmt_2262_branch_req_0); -- 
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_1786/ifx_xelse151_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_1786/ifx_xelse151_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1786/merge_stmt_2290_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1786/merge_stmt_2290_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_1786/merge_stmt_2290_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_1786/merge_stmt_2290_PhiAck/dummy
      -- CP-element group 85: 	 branch_block_stmt_1786/merge_stmt_2290__exit__
      -- CP-element group 85: 	 branch_block_stmt_1786/assign_stmt_2295__entry__
      -- CP-element group 85: 	 branch_block_stmt_1786/if_stmt_2262_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_1786/if_stmt_2262_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_1786/ifx_xelse151_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_1786/assign_stmt_2295/$entry
      -- CP-element group 85: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Sample/req
      -- 
    if_choice_transition_5567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2262_branch_ack_1, ack => zeropad3D_C_CP_4749_elements(85)); -- 
    req_5584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(85), ack => WPIPE_Block2_complete_2292_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	114 
    -- CP-element group 86: 	116 
    -- CP-element group 86: 	117 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2269/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1786/if_stmt_2262_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_1786/if_stmt_2262_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185
      -- 
    else_choice_transition_5571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2262_branch_ack_0, ack => zeropad3D_C_CP_4749_elements(86)); -- 
    cr_5813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(86), ack => type_cast_2279_inst_req_1); -- 
    cr_5836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(86), ack => type_cast_2287_inst_req_1); -- 
    rr_5831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(86), ack => type_cast_2287_inst_req_0); -- 
    rr_5808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(86), ack => type_cast_2279_inst_req_0); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Update/req
      -- 
    ack_5585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_complete_2292_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(87)); -- 
    req_5589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(87), ack => WPIPE_Block2_complete_2292_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1786/merge_stmt_2297_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1786/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_1786/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_1786/merge_stmt_2297_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1786/merge_stmt_2297_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_1786/merge_stmt_2297_PhiAck/dummy
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_1786/$exit
      -- CP-element group 88: 	 branch_block_stmt_1786/branch_block_stmt_1786__exit__
      -- CP-element group 88: 	 branch_block_stmt_1786/assign_stmt_2295__exit__
      -- CP-element group 88: 	 branch_block_stmt_1786/return__
      -- CP-element group 88: 	 branch_block_stmt_1786/merge_stmt_2297__exit__
      -- CP-element group 88: 	 branch_block_stmt_1786/assign_stmt_2295/$exit
      -- CP-element group 88: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1786/assign_stmt_2295/WPIPE_Block2_complete_2292_Update/ack
      -- 
    ack_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_complete_2292_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(88)); -- 
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	94 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1940/$exit
      -- CP-element group 89: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1944_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_req
      -- 
    phi_stmt_1940_req_5601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1940_req_5601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(89), ack => phi_stmt_1940_req_0); -- 
    -- Element group zeropad3D_C_CP_4749_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_4749_elements(32), ack => zeropad3D_C_CP_4749_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	32 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Sample/ra
      -- 
    ra_5618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/Update/ca
      -- 
    ca_5623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/$exit
      -- CP-element group 92: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/$exit
      -- CP-element group 92: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_req
      -- 
    phi_stmt_1934_req_5624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1934_req_5624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(92), ack => phi_stmt_1934_req_0); -- 
    zeropad3D_C_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(90) & zeropad3D_C_CP_4749_elements(91);
      gj_zeropad3D_C_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	32 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1927/$exit
      -- CP-element group 93: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1931_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_req
      -- 
    phi_stmt_1927_req_5632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1927_req_5632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(93), ack => phi_stmt_1927_req_0); -- 
    -- Element group zeropad3D_C_CP_4749_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_4749_elements(32), ack => zeropad3D_C_CP_4749_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	105 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1786/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(89) & zeropad3D_C_CP_4749_elements(92) & zeropad3D_C_CP_4749_elements(93);
      gj_zeropad3D_C_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Sample/ra
      -- 
    ra_5652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1946_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/Update/ca
      -- 
    ca_5657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1946_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/$exit
      -- CP-element group 97: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/$exit
      -- CP-element group 97: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_sources/type_cast_1946/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1940/phi_stmt_1940_req
      -- 
    phi_stmt_1940_req_5658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1940_req_5658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(97), ack => phi_stmt_1940_req_1); -- 
    zeropad3D_C_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(95) & zeropad3D_C_CP_4749_elements(96);
      gj_zeropad3D_C_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Sample/ra
      -- 
    ra_5675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1939_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/Update/ca
      -- 
    ca_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1939_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/$exit
      -- CP-element group 100: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/$exit
      -- CP-element group 100: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1939/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1934/phi_stmt_1934_req
      -- 
    phi_stmt_1934_req_5681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1934_req_5681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(100), ack => phi_stmt_1934_req_1); -- 
    zeropad3D_C_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(98) & zeropad3D_C_CP_4749_elements(99);
      gj_zeropad3D_C_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Sample/ra
      -- 
    ra_5698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/Update/ca
      -- 
    ca_5703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/$exit
      -- CP-element group 103: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/$exit
      -- CP-element group 103: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_sources/type_cast_1933/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/phi_stmt_1927/phi_stmt_1927_req
      -- 
    phi_stmt_1927_req_5704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1927_req_5704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(103), ack => phi_stmt_1927_req_1); -- 
    zeropad3D_C_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(101) & zeropad3D_C_CP_4749_elements(102);
      gj_zeropad3D_C_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1786/ifx_xend185_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(97) & zeropad3D_C_CP_4749_elements(100) & zeropad3D_C_CP_4749_elements(103);
      gj_zeropad3D_C_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  merge  fork  transition  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	94 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1786/merge_stmt_1926_PhiReqMerge
      -- CP-element group 105: 	 branch_block_stmt_1786/merge_stmt_1926_PhiAck/$entry
      -- 
    zeropad3D_C_CP_4749_elements(105) <= OrReduce(zeropad3D_C_CP_4749_elements(94) & zeropad3D_C_CP_4749_elements(104));
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1786/merge_stmt_1926_PhiAck/phi_stmt_1927_ack
      -- 
    phi_stmt_1927_ack_5709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1927_ack_0, ack => zeropad3D_C_CP_4749_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1786/merge_stmt_1926_PhiAck/phi_stmt_1934_ack
      -- 
    phi_stmt_1934_ack_5710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1934_ack_0, ack => zeropad3D_C_CP_4749_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1786/merge_stmt_1926_PhiAck/phi_stmt_1940_ack
      -- 
    phi_stmt_1940_ack_5711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1940_ack_0, ack => zeropad3D_C_CP_4749_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	34 
    -- CP-element group 109: 	33 
    -- CP-element group 109:  members (10) 
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/$entry
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1786/merge_stmt_1926__exit__
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977__entry__
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1786/assign_stmt_1952_to_assign_stmt_1977/type_cast_1951_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_1786/merge_stmt_1926_PhiAck/$exit
      -- 
    rr_5031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(109), ack => type_cast_1951_inst_req_0); -- 
    cr_5036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(109), ack => type_cast_1951_inst_req_1); -- 
    zeropad3D_C_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(106) & zeropad3D_C_CP_4749_elements(107) & zeropad3D_C_CP_4749_elements(108);
      gj_zeropad3D_C_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  merge  fork  transition  place  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	36 
    -- CP-element group 110: 	40 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	53 
    -- CP-element group 110: 	51 
    -- CP-element group 110: 	43 
    -- CP-element group 110: 	47 
    -- CP-element group 110: 	44 
    -- CP-element group 110: 	42 
    -- CP-element group 110: 	41 
    -- CP-element group 110:  members (33) 
      -- CP-element group 110: 	 branch_block_stmt_1786/merge_stmt_2021__exit__
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077__entry__
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2025_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2030_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/type_cast_2064_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_update_start
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/array_obj_ref_2070_final_index_sum_regn_Update/req
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/addr_of_2071_complete/req
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/word_access_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/word_access_complete/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/assign_stmt_2026_to_assign_stmt_2077/ptr_deref_2074_Update/word_access_complete/word_0/cr
      -- CP-element group 110: 	 branch_block_stmt_1786/merge_stmt_2021_PhiReqMerge
      -- CP-element group 110: 	 branch_block_stmt_1786/merge_stmt_2021_PhiAck/$entry
      -- CP-element group 110: 	 branch_block_stmt_1786/merge_stmt_2021_PhiAck/$exit
      -- CP-element group 110: 	 branch_block_stmt_1786/merge_stmt_2021_PhiAck/dummy
      -- 
    rr_5103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => type_cast_2025_inst_req_0); -- 
    cr_5108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => type_cast_2025_inst_req_1); -- 
    rr_5117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => type_cast_2030_inst_req_0); -- 
    cr_5122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => type_cast_2030_inst_req_1); -- 
    cr_5136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => type_cast_2064_inst_req_1); -- 
    req_5167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => array_obj_ref_2070_index_offset_req_1); -- 
    req_5182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => addr_of_2071_final_reg_req_1); -- 
    cr_5232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(110), ack => ptr_deref_2074_store_0_req_1); -- 
    zeropad3D_C_CP_4749_elements(110) <= OrReduce(zeropad3D_C_CP_4749_elements(36) & zeropad3D_C_CP_4749_elements(40));
    -- CP-element group 111:  merge  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	54 
    -- CP-element group 111: 	74 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	75 
    -- CP-element group 111: 	76 
    -- CP-element group 111:  members (13) 
      -- CP-element group 111: 	 branch_block_stmt_1786/merge_stmt_2186_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_1786/merge_stmt_2186_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_1786/merge_stmt_2186_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_1786/merge_stmt_2186_PhiAck/dummy
      -- CP-element group 111: 	 branch_block_stmt_1786/merge_stmt_2186__exit__
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204__entry__
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/$entry
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1786/assign_stmt_2191_to_assign_stmt_2204/type_cast_2190_Update/cr
      -- 
    rr_5481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(111), ack => type_cast_2190_inst_req_0); -- 
    cr_5486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(111), ack => type_cast_2190_inst_req_1); -- 
    zeropad3D_C_CP_4749_elements(111) <= OrReduce(zeropad3D_C_CP_4749_elements(54) & zeropad3D_C_CP_4749_elements(74));
    -- CP-element group 112:  transition  output  delay-element  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	119 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_req
      -- CP-element group 112: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2275_konst_delay_trans
      -- CP-element group 112: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$exit
      -- CP-element group 112: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2269/$exit
      -- 
    phi_stmt_2269_req_5792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2269_req_5792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(112), ack => phi_stmt_2269_req_1); -- 
    -- Element group zeropad3D_C_CP_4749_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_4749_elements(86), ack => zeropad3D_C_CP_4749_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Sample/$exit
      -- 
    ra_5809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	86 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/Update/$exit
      -- 
    ca_5814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	119 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_req
      -- CP-element group 115: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/$exit
      -- CP-element group 115: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/$exit
      -- CP-element group 115: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2279/SplitProtocol/$exit
      -- 
    phi_stmt_2276_req_5815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2276_req_5815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(115), ack => phi_stmt_2276_req_0); -- 
    zeropad3D_C_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(113) & zeropad3D_C_CP_4749_elements(114);
      gj_zeropad3D_C_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Sample/$exit
      -- 
    ra_5832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	86 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/Update/$exit
      -- 
    ca_5837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/$exit
      -- CP-element group 118: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/$exit
      -- CP-element group 118: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2287/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_req
      -- 
    phi_stmt_2282_req_5838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2282_req_5838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(118), ack => phi_stmt_2282_req_1); -- 
    zeropad3D_C_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(116) & zeropad3D_C_CP_4749_elements(117);
      gj_zeropad3D_C_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	112 
    -- CP-element group 119: 	115 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	130 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1786/ifx_xelse151_ifx_xend185_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(112) & zeropad3D_C_CP_4749_elements(115) & zeropad3D_C_CP_4749_elements(118);
      gj_zeropad3D_C_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/$exit
      -- 
    ra_5858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/ca
      -- 
    ca_5863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	129 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/$exit
      -- CP-element group 122: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/$exit
      -- CP-element group 122: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2269/phi_stmt_2269_req
      -- 
    phi_stmt_2269_req_5864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2269_req_5864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(122), ack => phi_stmt_2269_req_0); -- 
    zeropad3D_C_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(120) & zeropad3D_C_CP_4749_elements(121);
      gj_zeropad3D_C_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Sample/ra
      -- 
    ra_5881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2281_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/Update/ca
      -- 
    ca_5886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2281_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/$exit
      -- CP-element group 125: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/type_cast_2281/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_req
      -- CP-element group 125: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/phi_stmt_2276_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2276/$exit
      -- 
    phi_stmt_2276_req_5887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2276_req_5887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(125), ack => phi_stmt_2276_req_1); -- 
    zeropad3D_C_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(123) & zeropad3D_C_CP_4749_elements(124);
      gj_zeropad3D_C_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Sample/$exit
      -- 
    ra_5904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2285_inst_ack_0, ack => zeropad3D_C_CP_4749_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	77 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Update/ca
      -- CP-element group 127: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/Update/$exit
      -- 
    ca_5909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2285_inst_ack_1, ack => zeropad3D_C_CP_4749_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/$exit
      -- CP-element group 128: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_req
      -- CP-element group 128: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2285/$exit
      -- CP-element group 128: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$exit
      -- 
    phi_stmt_2282_req_5910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2282_req_5910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4749_elements(128), ack => phi_stmt_2282_req_0); -- 
    zeropad3D_C_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(126) & zeropad3D_C_CP_4749_elements(127);
      gj_zeropad3D_C_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1786/ifx_xthen146_ifx_xend185_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(122) & zeropad3D_C_CP_4749_elements(125) & zeropad3D_C_CP_4749_elements(128);
      gj_zeropad3D_C_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1786/merge_stmt_2268_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1786/merge_stmt_2268_PhiAck/$entry
      -- 
    zeropad3D_C_CP_4749_elements(130) <= OrReduce(zeropad3D_C_CP_4749_elements(119) & zeropad3D_C_CP_4749_elements(129));
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1786/merge_stmt_2268_PhiAck/phi_stmt_2269_ack
      -- 
    phi_stmt_2269_ack_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2269_ack_0, ack => zeropad3D_C_CP_4749_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1786/merge_stmt_2268_PhiAck/phi_stmt_2276_ack
      -- 
    phi_stmt_2276_ack_5916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2276_ack_0, ack => zeropad3D_C_CP_4749_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1786/merge_stmt_2268_PhiAck/phi_stmt_2282_ack
      -- 
    phi_stmt_2282_ack_5917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2282_ack_0, ack => zeropad3D_C_CP_4749_elements(133)); -- 
    -- CP-element group 134:  join  transition  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	1 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1786/merge_stmt_2268_PhiAck/$exit
      -- 
    zeropad3D_C_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4749_elements(131) & zeropad3D_C_CP_4749_elements(132) & zeropad3D_C_CP_4749_elements(133);
      gj_zeropad3D_C_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4749_elements(134), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1860_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1922_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2058_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2141_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2166_wire : std_logic_vector(31 downto 0);
    signal R_idxprom131_2152_resized : std_logic_vector(13 downto 0);
    signal R_idxprom131_2152_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom136_2177_resized : std_logic_vector(13 downto 0);
    signal R_idxprom136_2177_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2069_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2069_scaled : std_logic_vector(13 downto 0);
    signal add103_2109 : std_logic_vector(31 downto 0);
    signal add112_2114 : std_logic_vector(31 downto 0);
    signal add122_2129 : std_logic_vector(31 downto 0);
    signal add128_2134 : std_logic_vector(31 downto 0);
    signal add141_2197 : std_logic_vector(31 downto 0);
    signal add149_2217 : std_logic_vector(15 downto 0);
    signal add160_1879 : std_logic_vector(31 downto 0);
    signal add176_1894 : std_logic_vector(31 downto 0);
    signal add74_1904 : std_logic_vector(31 downto 0);
    signal add85_2046 : std_logic_vector(31 downto 0);
    signal add91_2051 : std_logic_vector(31 downto 0);
    signal add_1899 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2070_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2070_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2070_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2070_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2070_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2070_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2153_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2153_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2153_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2153_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2153_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2153_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_root_address : std_logic_vector(13 downto 0);
    signal arrayidx132_2155 : std_logic_vector(31 downto 0);
    signal arrayidx137_2180 : std_logic_vector(31 downto 0);
    signal arrayidx_2072 : std_logic_vector(31 downto 0);
    signal call1_1792 : std_logic_vector(7 downto 0);
    signal call2_1795 : std_logic_vector(7 downto 0);
    signal call3_1798 : std_logic_vector(7 downto 0);
    signal call4_1801 : std_logic_vector(7 downto 0);
    signal call5_1804 : std_logic_vector(7 downto 0);
    signal call6_1807 : std_logic_vector(7 downto 0);
    signal call_1789 : std_logic_vector(7 downto 0);
    signal cmp144_2204 : std_logic_vector(0 downto 0);
    signal cmp161_2235 : std_logic_vector(0 downto 0);
    signal cmp177_2261 : std_logic_vector(0 downto 0);
    signal cmp57_1972 : std_logic_vector(0 downto 0);
    signal cmp64_1996 : std_logic_vector(0 downto 0);
    signal cmp64x_xnot_2002 : std_logic_vector(0 downto 0);
    signal cmp75_2009 : std_logic_vector(0 downto 0);
    signal cmp_1959 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_1965 : std_logic_vector(0 downto 0);
    signal conv105_1924 : std_logic_vector(31 downto 0);
    signal conv140_2191 : std_logic_vector(31 downto 0);
    signal conv154_2230 : std_logic_vector(31 downto 0);
    signal conv169_2256 : std_logic_vector(31 downto 0);
    signal conv171_1883 : std_logic_vector(31 downto 0);
    signal conv31_1822 : std_logic_vector(31 downto 0);
    signal conv33_1826 : std_logic_vector(31 downto 0);
    signal conv37_1830 : std_logic_vector(31 downto 0);
    signal conv39_1834 : std_logic_vector(31 downto 0);
    signal conv46_1952 : std_logic_vector(31 downto 0);
    signal conv48_1843 : std_logic_vector(31 downto 0);
    signal conv61_1989 : std_logic_vector(31 downto 0);
    signal conv79_2026 : std_logic_vector(31 downto 0);
    signal conv81_1847 : std_logic_vector(31 downto 0);
    signal conv83_2031 : std_logic_vector(31 downto 0);
    signal conv87_1862 : std_logic_vector(31 downto 0);
    signal conv95_2084 : std_logic_vector(31 downto 0);
    signal conv_1812 : std_logic_vector(15 downto 0);
    signal div157_1868 : std_logic_vector(31 downto 0);
    signal div172_1889 : std_logic_vector(31 downto 0);
    signal div_1818 : std_logic_vector(15 downto 0);
    signal idxprom131_2148 : std_logic_vector(63 downto 0);
    signal idxprom136_2173 : std_logic_vector(63 downto 0);
    signal idxprom_2065 : std_logic_vector(63 downto 0);
    signal inc166_2239 : std_logic_vector(15 downto 0);
    signal inc166x_xix_x2_2244 : std_logic_vector(15 downto 0);
    signal inc_2225 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_2276 : std_logic_vector(15 downto 0);
    signal ix_x2_1934 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_2282 : std_logic_vector(15 downto 0);
    signal jx_x1_1940 : std_logic_vector(15 downto 0);
    signal jx_x2_2251 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_2269 : std_logic_vector(15 downto 0);
    signal kx_x1_1927 : std_logic_vector(15 downto 0);
    signal mul102_2094 : std_logic_vector(31 downto 0);
    signal mul111_2104 : std_logic_vector(31 downto 0);
    signal mul121_2119 : std_logic_vector(31 downto 0);
    signal mul127_2124 : std_logic_vector(31 downto 0);
    signal mul40_1839 : std_logic_vector(31 downto 0);
    signal mul84_2036 : std_logic_vector(31 downto 0);
    signal mul90_2041 : std_logic_vector(31 downto 0);
    signal mul_1910 : std_logic_vector(31 downto 0);
    signal orx_xcond191_2014 : std_logic_vector(0 downto 0);
    signal orx_xcond_1977 : std_logic_vector(0 downto 0);
    signal ptr_deref_2074_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2074_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2074_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2074_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2074_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2074_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2158_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2158_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2158_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2158_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2158_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2182_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2182_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext190_1853 : std_logic_vector(31 downto 0);
    signal sext_1915 : std_logic_vector(31 downto 0);
    signal shl_1874 : std_logic_vector(31 downto 0);
    signal shr130_2143 : std_logic_vector(31 downto 0);
    signal shr135_2168 : std_logic_vector(31 downto 0);
    signal shr_2060 : std_logic_vector(31 downto 0);
    signal sub110_2099 : std_logic_vector(31 downto 0);
    signal sub_2089 : std_logic_vector(31 downto 0);
    signal tmp133_2159 : std_logic_vector(63 downto 0);
    signal type_cast_1816_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1851_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1856_wire : std_logic_vector(31 downto 0);
    signal type_cast_1859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1866_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1872_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1887_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1908_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1918_wire : std_logic_vector(31 downto 0);
    signal type_cast_1921_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1931_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1933_wire : std_logic_vector(15 downto 0);
    signal type_cast_1937_wire : std_logic_vector(15 downto 0);
    signal type_cast_1939_wire : std_logic_vector(15 downto 0);
    signal type_cast_1944_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1946_wire : std_logic_vector(15 downto 0);
    signal type_cast_1950_wire : std_logic_vector(31 downto 0);
    signal type_cast_1955_wire : std_logic_vector(31 downto 0);
    signal type_cast_1957_wire : std_logic_vector(31 downto 0);
    signal type_cast_1963_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1968_wire : std_logic_vector(31 downto 0);
    signal type_cast_1970_wire : std_logic_vector(31 downto 0);
    signal type_cast_1987_wire : std_logic_vector(31 downto 0);
    signal type_cast_1992_wire : std_logic_vector(31 downto 0);
    signal type_cast_1994_wire : std_logic_vector(31 downto 0);
    signal type_cast_2000_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2005_wire : std_logic_vector(31 downto 0);
    signal type_cast_2007_wire : std_logic_vector(31 downto 0);
    signal type_cast_2024_wire : std_logic_vector(31 downto 0);
    signal type_cast_2029_wire : std_logic_vector(31 downto 0);
    signal type_cast_2054_wire : std_logic_vector(31 downto 0);
    signal type_cast_2057_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2063_wire : std_logic_vector(63 downto 0);
    signal type_cast_2076_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2082_wire : std_logic_vector(31 downto 0);
    signal type_cast_2137_wire : std_logic_vector(31 downto 0);
    signal type_cast_2140_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2146_wire : std_logic_vector(63 downto 0);
    signal type_cast_2162_wire : std_logic_vector(31 downto 0);
    signal type_cast_2165_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2171_wire : std_logic_vector(63 downto 0);
    signal type_cast_2189_wire : std_logic_vector(31 downto 0);
    signal type_cast_2195_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2200_wire : std_logic_vector(31 downto 0);
    signal type_cast_2202_wire : std_logic_vector(31 downto 0);
    signal type_cast_2215_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2223_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2228_wire : std_logic_vector(31 downto 0);
    signal type_cast_2248_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2254_wire : std_logic_vector(31 downto 0);
    signal type_cast_2272_wire : std_logic_vector(15 downto 0);
    signal type_cast_2275_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2279_wire : std_logic_vector(15 downto 0);
    signal type_cast_2281_wire : std_logic_vector(15 downto 0);
    signal type_cast_2285_wire : std_logic_vector(15 downto 0);
    signal type_cast_2287_wire : std_logic_vector(15 downto 0);
    signal type_cast_2294_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_2070_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2070_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2070_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2070_resized_base_address <= "00000000000000";
    array_obj_ref_2153_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2153_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2153_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2153_resized_base_address <= "00000000000000";
    array_obj_ref_2178_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2178_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2178_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2178_resized_base_address <= "00000000000000";
    ptr_deref_2074_word_offset_0 <= "00000000000000";
    ptr_deref_2158_word_offset_0 <= "00000000000000";
    ptr_deref_2182_word_offset_0 <= "00000000000000";
    type_cast_1816_wire_constant <= "0000000000000010";
    type_cast_1851_wire_constant <= "00000000000000000000000000010000";
    type_cast_1859_wire_constant <= "00000000000000000000000000010000";
    type_cast_1866_wire_constant <= "00000000000000000000000000000001";
    type_cast_1872_wire_constant <= "00000000000000000000000000000001";
    type_cast_1887_wire_constant <= "00000000000000000000000000000001";
    type_cast_1908_wire_constant <= "00000000000000000000000000010000";
    type_cast_1921_wire_constant <= "00000000000000000000000000010000";
    type_cast_1931_wire_constant <= "0000000000000000";
    type_cast_1944_wire_constant <= "0000000000000000";
    type_cast_1963_wire_constant <= "1";
    type_cast_2000_wire_constant <= "1";
    type_cast_2057_wire_constant <= "00000000000000000000000000000010";
    type_cast_2076_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2140_wire_constant <= "00000000000000000000000000000010";
    type_cast_2165_wire_constant <= "00000000000000000000000000000010";
    type_cast_2195_wire_constant <= "00000000000000000000000000000100";
    type_cast_2215_wire_constant <= "0000000000000100";
    type_cast_2223_wire_constant <= "0000000000000001";
    type_cast_2248_wire_constant <= "0000000000000000";
    type_cast_2275_wire_constant <= "0000000000000000";
    type_cast_2294_wire_constant <= "00000001";
    phi_stmt_1927: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1931_wire_constant & type_cast_1933_wire;
      req <= phi_stmt_1927_req_0 & phi_stmt_1927_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1927",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1927_ack_0,
          idata => idata,
          odata => kx_x1_1927,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1927
    phi_stmt_1934: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1937_wire & type_cast_1939_wire;
      req <= phi_stmt_1934_req_0 & phi_stmt_1934_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1934",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1934_ack_0,
          idata => idata,
          odata => ix_x2_1934,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1934
    phi_stmt_1940: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1944_wire_constant & type_cast_1946_wire;
      req <= phi_stmt_1940_req_0 & phi_stmt_1940_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1940",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1940_ack_0,
          idata => idata,
          odata => jx_x1_1940,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1940
    phi_stmt_2269: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2272_wire & type_cast_2275_wire_constant;
      req <= phi_stmt_2269_req_0 & phi_stmt_2269_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2269",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2269_ack_0,
          idata => idata,
          odata => kx_x0x_xph_2269,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2269
    phi_stmt_2276: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2279_wire & type_cast_2281_wire;
      req <= phi_stmt_2276_req_0 & phi_stmt_2276_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2276",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2276_ack_0,
          idata => idata,
          odata => ix_x1x_xph_2276,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2276
    phi_stmt_2282: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2285_wire & type_cast_2287_wire;
      req <= phi_stmt_2282_req_0 & phi_stmt_2282_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2282",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2282_ack_0,
          idata => idata,
          odata => jx_x0x_xph_2282,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2282
    -- flow-through select operator MUX_2250_inst
    jx_x2_2251 <= type_cast_2248_wire_constant when (cmp161_2235(0) /=  '0') else inc_2225;
    addr_of_2071_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2071_final_reg_req_0;
      addr_of_2071_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2071_final_reg_req_1;
      addr_of_2071_final_reg_ack_1<= rack(0);
      addr_of_2071_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2071_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2070_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2072,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2154_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2154_final_reg_req_0;
      addr_of_2154_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2154_final_reg_req_1;
      addr_of_2154_final_reg_ack_1<= rack(0);
      addr_of_2154_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2154_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2153_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx132_2155,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2179_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2179_final_reg_req_0;
      addr_of_2179_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2179_final_reg_req_1;
      addr_of_2179_final_reg_ack_1<= rack(0);
      addr_of_2179_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2179_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2178_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx137_2180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1811_inst_req_0;
      type_cast_1811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1811_inst_req_1;
      type_cast_1811_inst_ack_1<= rack(0);
      type_cast_1811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1812,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1821_inst_req_0;
      type_cast_1821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1821_inst_req_1;
      type_cast_1821_inst_ack_1<= rack(0);
      type_cast_1821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_1822,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1825_inst_req_0;
      type_cast_1825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1825_inst_req_1;
      type_cast_1825_inst_ack_1<= rack(0);
      type_cast_1825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1829_inst_req_0;
      type_cast_1829_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1829_inst_req_1;
      type_cast_1829_inst_ack_1<= rack(0);
      type_cast_1829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1829_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_1830,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1833_inst_req_0;
      type_cast_1833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1833_inst_req_1;
      type_cast_1833_inst_ack_1<= rack(0);
      type_cast_1833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_1801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1842_inst_req_0;
      type_cast_1842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1842_inst_req_1;
      type_cast_1842_inst_ack_1<= rack(0);
      type_cast_1842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_1843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1846_inst_req_0;
      type_cast_1846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1846_inst_req_1;
      type_cast_1846_inst_ack_1<= rack(0);
      type_cast_1846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1847,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1856_inst
    process(sext190_1853) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext190_1853(31 downto 0);
      type_cast_1856_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1861_inst
    process(ASHR_i32_i32_1860_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1860_wire(31 downto 0);
      conv87_1862 <= tmp_var; -- 
    end process;
    type_cast_1882_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1882_inst_req_0;
      type_cast_1882_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1882_inst_req_1;
      type_cast_1882_inst_ack_1<= rack(0);
      type_cast_1882_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1882_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_1883,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1918_inst
    process(sext_1915) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1915(31 downto 0);
      type_cast_1918_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1923_inst
    process(ASHR_i32_i32_1922_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1922_wire(31 downto 0);
      conv105_1924 <= tmp_var; -- 
    end process;
    type_cast_1933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1933_inst_req_0;
      type_cast_1933_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1933_inst_req_1;
      type_cast_1933_inst_ack_1<= rack(0);
      type_cast_1933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_2269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1933_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1937_inst_req_0;
      type_cast_1937_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1937_inst_req_1;
      type_cast_1937_inst_ack_1<= rack(0);
      type_cast_1937_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1937_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1818,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1937_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1939_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1939_inst_req_0;
      type_cast_1939_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1939_inst_req_1;
      type_cast_1939_inst_ack_1<= rack(0);
      type_cast_1939_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1939_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_2276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1939_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1946_inst_req_0;
      type_cast_1946_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1946_inst_req_1;
      type_cast_1946_inst_ack_1<= rack(0);
      type_cast_1946_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1946_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_2282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1946_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1951_inst_req_0;
      type_cast_1951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1951_inst_req_1;
      type_cast_1951_inst_ack_1<= rack(0);
      type_cast_1951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1950_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_1952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1955_inst
    process(conv46_1952) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_1952(31 downto 0);
      type_cast_1955_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1957_inst
    process(conv48_1843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_1843(31 downto 0);
      type_cast_1957_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1968_inst
    process(conv46_1952) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_1952(31 downto 0);
      type_cast_1968_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1970_inst
    process(add_1899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_1899(31 downto 0);
      type_cast_1970_wire <= tmp_var; -- 
    end process;
    type_cast_1988_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1988_inst_req_0;
      type_cast_1988_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1988_inst_req_1;
      type_cast_1988_inst_ack_1<= rack(0);
      type_cast_1988_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1988_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1987_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1989,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1992_inst
    process(conv61_1989) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv61_1989(31 downto 0);
      type_cast_1992_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1994_inst
    process(conv48_1843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_1843(31 downto 0);
      type_cast_1994_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2005_inst
    process(conv61_1989) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv61_1989(31 downto 0);
      type_cast_2005_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2007_inst
    process(add74_1904) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add74_1904(31 downto 0);
      type_cast_2007_wire <= tmp_var; -- 
    end process;
    type_cast_2025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2025_inst_req_0;
      type_cast_2025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2025_inst_req_1;
      type_cast_2025_inst_ack_1<= rack(0);
      type_cast_2025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2024_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_2026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2030_inst_req_0;
      type_cast_2030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2030_inst_req_1;
      type_cast_2030_inst_ack_1<= rack(0);
      type_cast_2030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2029_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_2031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2054_inst
    process(add91_2051) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add91_2051(31 downto 0);
      type_cast_2054_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2059_inst
    process(ASHR_i32_i32_2058_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2058_wire(31 downto 0);
      shr_2060 <= tmp_var; -- 
    end process;
    type_cast_2064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2064_inst_req_0;
      type_cast_2064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2064_inst_req_1;
      type_cast_2064_inst_ack_1<= rack(0);
      type_cast_2064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2063_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2083_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2083_inst_req_0;
      type_cast_2083_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2083_inst_req_1;
      type_cast_2083_inst_ack_1<= rack(0);
      type_cast_2083_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2083_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2082_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2137_inst
    process(add112_2114) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add112_2114(31 downto 0);
      type_cast_2137_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2142_inst
    process(ASHR_i32_i32_2141_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2141_wire(31 downto 0);
      shr130_2143 <= tmp_var; -- 
    end process;
    type_cast_2147_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2147_inst_req_0;
      type_cast_2147_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2147_inst_req_1;
      type_cast_2147_inst_ack_1<= rack(0);
      type_cast_2147_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2147_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2146_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom131_2148,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2162_inst
    process(add128_2134) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add128_2134(31 downto 0);
      type_cast_2162_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2167_inst
    process(ASHR_i32_i32_2166_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2166_wire(31 downto 0);
      shr135_2168 <= tmp_var; -- 
    end process;
    type_cast_2172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2172_inst_req_0;
      type_cast_2172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2172_inst_req_1;
      type_cast_2172_inst_ack_1<= rack(0);
      type_cast_2172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2171_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom136_2173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2190_inst_req_0;
      type_cast_2190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2190_inst_req_1;
      type_cast_2190_inst_ack_1<= rack(0);
      type_cast_2190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2189_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_2191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2200_inst
    process(add141_2197) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add141_2197(31 downto 0);
      type_cast_2200_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2202_inst
    process(conv31_1822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv31_1822(31 downto 0);
      type_cast_2202_wire <= tmp_var; -- 
    end process;
    type_cast_2229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2229_inst_req_0;
      type_cast_2229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2229_inst_req_1;
      type_cast_2229_inst_ack_1<= rack(0);
      type_cast_2229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2228_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_2230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2238_inst_req_0;
      type_cast_2238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2238_inst_req_1;
      type_cast_2238_inst_ack_1<= rack(0);
      type_cast_2238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp161_2235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc166_2239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2255_inst_req_0;
      type_cast_2255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2255_inst_req_1;
      type_cast_2255_inst_ack_1<= rack(0);
      type_cast_2255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2254_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv169_2256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2272_inst_req_0;
      type_cast_2272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2272_inst_req_1;
      type_cast_2272_inst_ack_1<= rack(0);
      type_cast_2272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add149_2217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2272_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2279_inst_req_0;
      type_cast_2279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2279_inst_req_1;
      type_cast_2279_inst_ack_1<= rack(0);
      type_cast_2279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc166x_xix_x2_2244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2279_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2281_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2281_inst_req_0;
      type_cast_2281_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2281_inst_req_1;
      type_cast_2281_inst_ack_1<= rack(0);
      type_cast_2281_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2281_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_1934,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2281_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2285_inst_req_0;
      type_cast_2285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2285_inst_req_1;
      type_cast_2285_inst_ack_1<= rack(0);
      type_cast_2285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_1940,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2285_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2287_inst_req_0;
      type_cast_2287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2287_inst_req_1;
      type_cast_2287_inst_ack_1<= rack(0);
      type_cast_2287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_2251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2287_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2070_index_1_rename
    process(R_idxprom_2069_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2069_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2069_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2070_index_1_resize
    process(idxprom_2065) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2065;
      ov := iv(13 downto 0);
      R_idxprom_2069_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2070_root_address_inst
    process(array_obj_ref_2070_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2070_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2070_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2153_index_1_rename
    process(R_idxprom131_2152_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom131_2152_resized;
      ov(13 downto 0) := iv;
      R_idxprom131_2152_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2153_index_1_resize
    process(idxprom131_2148) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom131_2148;
      ov := iv(13 downto 0);
      R_idxprom131_2152_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2153_root_address_inst
    process(array_obj_ref_2153_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2153_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2153_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2178_index_1_rename
    process(R_idxprom136_2177_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom136_2177_resized;
      ov(13 downto 0) := iv;
      R_idxprom136_2177_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2178_index_1_resize
    process(idxprom136_2173) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom136_2173;
      ov := iv(13 downto 0);
      R_idxprom136_2177_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2178_root_address_inst
    process(array_obj_ref_2178_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2178_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2178_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2074_addr_0
    process(ptr_deref_2074_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2074_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2074_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2074_base_resize
    process(arrayidx_2072) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2072;
      ov := iv(13 downto 0);
      ptr_deref_2074_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2074_gather_scatter
    process(type_cast_2076_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2076_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2074_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2074_root_address_inst
    process(ptr_deref_2074_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2074_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2074_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2158_addr_0
    process(ptr_deref_2158_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2158_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2158_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2158_base_resize
    process(arrayidx132_2155) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx132_2155;
      ov := iv(13 downto 0);
      ptr_deref_2158_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2158_gather_scatter
    process(ptr_deref_2158_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2158_data_0;
      ov(63 downto 0) := iv;
      tmp133_2159 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2158_root_address_inst
    process(ptr_deref_2158_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2158_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2158_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_addr_0
    process(ptr_deref_2182_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2182_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2182_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_base_resize
    process(arrayidx137_2180) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx137_2180;
      ov := iv(13 downto 0);
      ptr_deref_2182_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_gather_scatter
    process(tmp133_2159) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp133_2159;
      ov(63 downto 0) := iv;
      ptr_deref_2182_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_root_address_inst
    process(ptr_deref_2182_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2182_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2182_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1978_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_1977;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1978_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1978_branch_req_0,
          ack0 => if_stmt_1978_branch_ack_0,
          ack1 => if_stmt_1978_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2015_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond191_2014;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2015_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2015_branch_req_0,
          ack0 => if_stmt_2015_branch_ack_0,
          ack1 => if_stmt_2015_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2205_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp144_2204;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2205_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2205_branch_req_0,
          ack0 => if_stmt_2205_branch_ack_0,
          ack1 => if_stmt_2205_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2262_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp177_2261;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2262_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2262_branch_req_0,
          ack0 => if_stmt_2262_branch_ack_0,
          ack1 => if_stmt_2262_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2216_inst
    process(kx_x1_1927) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_1927, type_cast_2215_wire_constant, tmp_var);
      add149_2217 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2224_inst
    process(jx_x1_1940) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_1940, type_cast_2223_wire_constant, tmp_var);
      inc_2225 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2243_inst
    process(inc166_2239, ix_x2_1934) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc166_2239, ix_x2_1934, tmp_var);
      inc166x_xix_x2_2244 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1878_inst
    process(shl_1874, div157_1868) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1874, div157_1868, tmp_var);
      add160_1879 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1893_inst
    process(shl_1874, div172_1889) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1874, div172_1889, tmp_var);
      add176_1894 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1898_inst
    process(conv48_1843, div172_1889) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv48_1843, div172_1889, tmp_var);
      add_1899 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1903_inst
    process(conv48_1843, div157_1868) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv48_1843, div157_1868, tmp_var);
      add74_1904 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2045_inst
    process(mul90_2041, conv79_2026) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul90_2041, conv79_2026, tmp_var);
      add85_2046 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2050_inst
    process(add85_2046, mul84_2036) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add85_2046, mul84_2036, tmp_var);
      add91_2051 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2108_inst
    process(mul111_2104, conv95_2084) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul111_2104, conv95_2084, tmp_var);
      add103_2109 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2113_inst
    process(add103_2109, mul102_2094) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add103_2109, mul102_2094, tmp_var);
      add112_2114 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2128_inst
    process(mul127_2124, conv95_2084) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul127_2124, conv95_2084, tmp_var);
      add122_2129 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2133_inst
    process(add122_2129, mul121_2119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add122_2129, mul121_2119, tmp_var);
      add128_2134 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2196_inst
    process(conv140_2191) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv140_2191, type_cast_2195_wire_constant, tmp_var);
      add141_2197 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1976_inst
    process(cmpx_xnot_1965, cmp57_1972) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_1965, cmp57_1972, tmp_var);
      orx_xcond_1977 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2013_inst
    process(cmp64x_xnot_2002, cmp75_2009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp64x_xnot_2002, cmp75_2009, tmp_var);
      orx_xcond191_2014 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1860_inst
    process(type_cast_1856_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1856_wire, type_cast_1859_wire_constant, tmp_var);
      ASHR_i32_i32_1860_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1922_inst
    process(type_cast_1918_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1918_wire, type_cast_1921_wire_constant, tmp_var);
      ASHR_i32_i32_1922_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2058_inst
    process(type_cast_2054_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2054_wire, type_cast_2057_wire_constant, tmp_var);
      ASHR_i32_i32_2058_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2141_inst
    process(type_cast_2137_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2137_wire, type_cast_2140_wire_constant, tmp_var);
      ASHR_i32_i32_2141_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2166_inst
    process(type_cast_2162_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2162_wire, type_cast_2165_wire_constant, tmp_var);
      ASHR_i32_i32_2166_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2234_inst
    process(conv154_2230, add160_1879) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv154_2230, add160_1879, tmp_var);
      cmp161_2235 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2260_inst
    process(conv169_2256, add176_1894) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv169_2256, add176_1894, tmp_var);
      cmp177_2261 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1817_inst
    process(conv_1812) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_1812, type_cast_1816_wire_constant, tmp_var);
      div_1818 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1867_inst
    process(conv33_1826) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv33_1826, type_cast_1866_wire_constant, tmp_var);
      div157_1868 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1888_inst
    process(conv171_1883) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv171_1883, type_cast_1887_wire_constant, tmp_var);
      div172_1889 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1838_inst
    process(conv37_1830, conv39_1834) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_1830, conv39_1834, tmp_var);
      mul40_1839 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1914_inst
    process(mul_1910, conv31_1822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1910, conv31_1822, tmp_var);
      sext_1915 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2035_inst
    process(conv83_2031, conv81_1847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv83_2031, conv81_1847, tmp_var);
      mul84_2036 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2040_inst
    process(conv46_1952, conv87_1862) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_1952, conv87_1862, tmp_var);
      mul90_2041 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2093_inst
    process(sub_2089, conv31_1822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_2089, conv31_1822, tmp_var);
      mul102_2094 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2103_inst
    process(sub110_2099, conv105_1924) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub110_2099, conv105_1924, tmp_var);
      mul111_2104 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2118_inst
    process(conv61_1989, conv81_1847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv61_1989, conv81_1847, tmp_var);
      mul121_2119 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2123_inst
    process(conv46_1952, conv87_1862) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_1952, conv87_1862, tmp_var);
      mul127_2124 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1852_inst
    process(mul40_1839) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul40_1839, type_cast_1851_wire_constant, tmp_var);
      sext190_1853 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1873_inst
    process(conv48_1843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_1843, type_cast_1872_wire_constant, tmp_var);
      shl_1874 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1909_inst
    process(conv33_1826) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv33_1826, type_cast_1908_wire_constant, tmp_var);
      mul_1910 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1958_inst
    process(type_cast_1955_wire, type_cast_1957_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1955_wire, type_cast_1957_wire, tmp_var);
      cmp_1959 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1971_inst
    process(type_cast_1968_wire, type_cast_1970_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1968_wire, type_cast_1970_wire, tmp_var);
      cmp57_1972 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1995_inst
    process(type_cast_1992_wire, type_cast_1994_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1992_wire, type_cast_1994_wire, tmp_var);
      cmp64_1996 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2008_inst
    process(type_cast_2005_wire, type_cast_2007_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2005_wire, type_cast_2007_wire, tmp_var);
      cmp75_2009 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2203_inst
    process(type_cast_2200_wire, type_cast_2202_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2200_wire, type_cast_2202_wire, tmp_var);
      cmp144_2204 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2088_inst
    process(conv61_1989, conv48_1843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv61_1989, conv48_1843, tmp_var);
      sub_2089 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2098_inst
    process(conv46_1952, conv48_1843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv46_1952, conv48_1843, tmp_var);
      sub110_2099 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1964_inst
    process(cmp_1959) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_1959, type_cast_1963_wire_constant, tmp_var);
      cmpx_xnot_1965 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2001_inst
    process(cmp64_1996) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp64_1996, type_cast_2000_wire_constant, tmp_var);
      cmp64x_xnot_2002 <= tmp_var; --
    end process;
    -- shared split operator group (46) : array_obj_ref_2070_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2069_scaled;
      array_obj_ref_2070_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2070_index_offset_req_0;
      array_obj_ref_2070_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2070_index_offset_req_1;
      array_obj_ref_2070_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_2153_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom131_2152_scaled;
      array_obj_ref_2153_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2153_index_offset_req_0;
      array_obj_ref_2153_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2153_index_offset_req_1;
      array_obj_ref_2153_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_2178_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom136_2177_scaled;
      array_obj_ref_2178_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2178_index_offset_req_0;
      array_obj_ref_2178_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2178_index_offset_req_1;
      array_obj_ref_2178_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- unary operator type_cast_1950_inst
    process(ix_x2_1934) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_1934, tmp_var);
      type_cast_1950_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1987_inst
    process(jx_x1_1940) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1940, tmp_var);
      type_cast_1987_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2024_inst
    process(kx_x1_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1927, tmp_var);
      type_cast_2024_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2029_inst
    process(jx_x1_1940) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1940, tmp_var);
      type_cast_2029_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2063_inst
    process(shr_2060) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2060, tmp_var);
      type_cast_2063_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2082_inst
    process(kx_x1_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1927, tmp_var);
      type_cast_2082_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2146_inst
    process(shr130_2143) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr130_2143, tmp_var);
      type_cast_2146_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2171_inst
    process(shr135_2168) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr135_2168, tmp_var);
      type_cast_2171_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2189_inst
    process(kx_x1_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1927, tmp_var);
      type_cast_2189_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2228_inst
    process(inc_2225) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2225, tmp_var);
      type_cast_2228_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2254_inst
    process(inc166x_xix_x2_2244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc166x_xix_x2_2244, tmp_var);
      type_cast_2254_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2158_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2158_load_0_req_0;
      ptr_deref_2158_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2158_load_0_req_1;
      ptr_deref_2158_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2158_word_address_0;
      ptr_deref_2158_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2074_store_0 ptr_deref_2182_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2074_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2182_store_0_req_0;
      ptr_deref_2074_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2182_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2074_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2182_store_0_req_1;
      ptr_deref_2074_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2182_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2074_word_address_0 & ptr_deref_2182_word_address_0;
      data_in <= ptr_deref_2074_data_0 & ptr_deref_2182_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_starting_1797_inst RPIPE_Block2_starting_1794_inst RPIPE_Block2_starting_1806_inst RPIPE_Block2_starting_1788_inst RPIPE_Block2_starting_1800_inst RPIPE_Block2_starting_1791_inst RPIPE_Block2_starting_1803_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block2_starting_1797_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_starting_1794_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_starting_1806_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_starting_1788_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_starting_1800_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_starting_1791_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_starting_1803_inst_req_0;
      RPIPE_Block2_starting_1797_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_starting_1794_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_starting_1806_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_starting_1788_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_starting_1800_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_starting_1791_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_starting_1803_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block2_starting_1797_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_starting_1794_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_starting_1806_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_starting_1788_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_starting_1800_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_starting_1791_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_starting_1803_inst_req_1;
      RPIPE_Block2_starting_1797_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_starting_1794_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_starting_1806_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_starting_1788_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_starting_1800_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_starting_1791_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_starting_1803_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call3_1798 <= data_out(55 downto 48);
      call2_1795 <= data_out(47 downto 40);
      call6_1807 <= data_out(39 downto 32);
      call_1789 <= data_out(31 downto 24);
      call4_1801 <= data_out(23 downto 16);
      call1_1792 <= data_out(15 downto 8);
      call5_1804 <= data_out(7 downto 0);
      Block2_starting_read_0_gI: SplitGuardInterface generic map(name => "Block2_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block2_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_starting_pipe_read_req(0),
          oack => Block2_starting_pipe_read_ack(0),
          odata => Block2_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_complete_2292_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_complete_2292_inst_req_0;
      WPIPE_Block2_complete_2292_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_complete_2292_inst_req_1;
      WPIPE_Block2_complete_2292_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2294_wire_constant;
      Block2_complete_write_0_gI: SplitGuardInterface generic map(name => "Block2_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_complete_pipe_write_req(0),
          oack => Block2_complete_pipe_write_ack(0),
          odata => Block2_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_C_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block3_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block3_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_D;
architecture zeropad3D_D_arch of zeropad3D_D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_D_CP_5934_start: Boolean;
  signal zeropad3D_D_CP_5934_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_2446_req_1 : boolean;
  signal type_cast_2747_inst_req_0 : boolean;
  signal type_cast_2708_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2303_inst_ack_0 : boolean;
  signal WPIPE_Block3_complete_2809_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2309_inst_ack_0 : boolean;
  signal type_cast_2690_inst_ack_1 : boolean;
  signal if_stmt_2779_branch_req_0 : boolean;
  signal type_cast_2708_inst_ack_1 : boolean;
  signal ptr_deref_2676_load_0_ack_0 : boolean;
  signal type_cast_2747_inst_ack_0 : boolean;
  signal type_cast_2756_inst_ack_1 : boolean;
  signal if_stmt_2779_branch_ack_1 : boolean;
  signal type_cast_2756_inst_req_1 : boolean;
  signal type_cast_2708_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2303_inst_ack_1 : boolean;
  signal RPIPE_Block3_starting_2303_inst_req_1 : boolean;
  signal type_cast_2756_inst_req_0 : boolean;
  signal addr_of_2697_final_reg_req_1 : boolean;
  signal RPIPE_Block3_starting_2318_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2318_inst_ack_1 : boolean;
  signal RPIPE_Block3_starting_2309_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2309_inst_ack_1 : boolean;
  signal addr_of_2697_final_reg_ack_0 : boolean;
  signal RPIPE_Block3_starting_2309_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2315_inst_ack_0 : boolean;
  signal addr_of_2697_final_reg_req_0 : boolean;
  signal RPIPE_Block3_starting_2312_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2312_inst_ack_1 : boolean;
  signal addr_of_2697_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_complete_2809_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2303_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2318_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2318_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2315_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2306_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2312_inst_ack_0 : boolean;
  signal type_cast_2690_inst_ack_0 : boolean;
  signal ptr_deref_2676_load_0_req_0 : boolean;
  signal WPIPE_Block3_complete_2809_inst_req_0 : boolean;
  signal type_cast_2690_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2315_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2315_inst_ack_1 : boolean;
  signal RPIPE_Block3_starting_2306_inst_req_0 : boolean;
  signal type_cast_2708_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2306_inst_ack_1 : boolean;
  signal type_cast_2756_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2312_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2306_inst_req_1 : boolean;
  signal WPIPE_Block3_complete_2809_inst_ack_1 : boolean;
  signal type_cast_2690_inst_req_0 : boolean;
  signal type_cast_2747_inst_req_1 : boolean;
  signal type_cast_2458_inst_req_0 : boolean;
  signal type_cast_2458_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2321_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2321_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2321_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2321_inst_ack_1 : boolean;
  signal if_stmt_2779_branch_ack_0 : boolean;
  signal type_cast_2326_inst_req_0 : boolean;
  signal ptr_deref_2700_store_0_ack_1 : boolean;
  signal type_cast_2326_inst_ack_0 : boolean;
  signal type_cast_2326_inst_req_1 : boolean;
  signal ptr_deref_2700_store_0_req_1 : boolean;
  signal type_cast_2326_inst_ack_1 : boolean;
  signal array_obj_ref_2696_index_offset_ack_1 : boolean;
  signal type_cast_2747_inst_ack_1 : boolean;
  signal type_cast_2336_inst_req_0 : boolean;
  signal type_cast_2336_inst_ack_0 : boolean;
  signal type_cast_2336_inst_req_1 : boolean;
  signal type_cast_2336_inst_ack_1 : boolean;
  signal if_stmt_2723_branch_ack_0 : boolean;
  signal array_obj_ref_2696_index_offset_req_1 : boolean;
  signal type_cast_2772_inst_ack_1 : boolean;
  signal type_cast_2346_inst_req_0 : boolean;
  signal type_cast_2346_inst_ack_0 : boolean;
  signal type_cast_2772_inst_req_1 : boolean;
  signal type_cast_2346_inst_req_1 : boolean;
  signal type_cast_2346_inst_ack_1 : boolean;
  signal if_stmt_2723_branch_ack_1 : boolean;
  signal array_obj_ref_2696_index_offset_ack_0 : boolean;
  signal array_obj_ref_2696_index_offset_req_0 : boolean;
  signal type_cast_2350_inst_req_0 : boolean;
  signal type_cast_2350_inst_ack_0 : boolean;
  signal type_cast_2350_inst_req_1 : boolean;
  signal type_cast_2350_inst_ack_1 : boolean;
  signal ptr_deref_2676_load_0_ack_1 : boolean;
  signal type_cast_2772_inst_ack_0 : boolean;
  signal type_cast_2354_inst_req_0 : boolean;
  signal ptr_deref_2700_store_0_ack_0 : boolean;
  signal type_cast_2354_inst_ack_0 : boolean;
  signal type_cast_2772_inst_req_0 : boolean;
  signal type_cast_2354_inst_req_1 : boolean;
  signal ptr_deref_2700_store_0_req_0 : boolean;
  signal type_cast_2354_inst_ack_1 : boolean;
  signal ptr_deref_2676_load_0_req_1 : boolean;
  signal if_stmt_2723_branch_req_0 : boolean;
  signal type_cast_2358_inst_req_0 : boolean;
  signal type_cast_2358_inst_ack_0 : boolean;
  signal type_cast_2358_inst_req_1 : boolean;
  signal type_cast_2358_inst_ack_1 : boolean;
  signal type_cast_2367_inst_req_0 : boolean;
  signal type_cast_2367_inst_ack_0 : boolean;
  signal type_cast_2367_inst_req_1 : boolean;
  signal type_cast_2367_inst_ack_1 : boolean;
  signal type_cast_2371_inst_req_0 : boolean;
  signal type_cast_2371_inst_ack_0 : boolean;
  signal type_cast_2371_inst_req_1 : boolean;
  signal type_cast_2371_inst_ack_1 : boolean;
  signal type_cast_2401_inst_req_0 : boolean;
  signal type_cast_2401_inst_ack_0 : boolean;
  signal type_cast_2401_inst_req_1 : boolean;
  signal type_cast_2401_inst_ack_1 : boolean;
  signal type_cast_2469_inst_req_0 : boolean;
  signal type_cast_2469_inst_ack_0 : boolean;
  signal type_cast_2469_inst_req_1 : boolean;
  signal type_cast_2469_inst_ack_1 : boolean;
  signal if_stmt_2496_branch_req_0 : boolean;
  signal if_stmt_2496_branch_ack_1 : boolean;
  signal if_stmt_2496_branch_ack_0 : boolean;
  signal type_cast_2506_inst_req_0 : boolean;
  signal type_cast_2506_inst_ack_0 : boolean;
  signal type_cast_2506_inst_req_1 : boolean;
  signal type_cast_2506_inst_ack_1 : boolean;
  signal if_stmt_2533_branch_req_0 : boolean;
  signal if_stmt_2533_branch_ack_1 : boolean;
  signal if_stmt_2533_branch_ack_0 : boolean;
  signal type_cast_2543_inst_req_0 : boolean;
  signal type_cast_2543_inst_ack_0 : boolean;
  signal type_cast_2543_inst_req_1 : boolean;
  signal type_cast_2543_inst_ack_1 : boolean;
  signal type_cast_2548_inst_req_0 : boolean;
  signal type_cast_2548_inst_ack_0 : boolean;
  signal type_cast_2548_inst_req_1 : boolean;
  signal type_cast_2548_inst_ack_1 : boolean;
  signal type_cast_2582_inst_req_0 : boolean;
  signal type_cast_2582_inst_ack_0 : boolean;
  signal type_cast_2582_inst_req_1 : boolean;
  signal type_cast_2582_inst_ack_1 : boolean;
  signal array_obj_ref_2588_index_offset_req_0 : boolean;
  signal array_obj_ref_2588_index_offset_ack_0 : boolean;
  signal array_obj_ref_2588_index_offset_req_1 : boolean;
  signal array_obj_ref_2588_index_offset_ack_1 : boolean;
  signal addr_of_2589_final_reg_req_0 : boolean;
  signal addr_of_2589_final_reg_ack_0 : boolean;
  signal addr_of_2589_final_reg_req_1 : boolean;
  signal addr_of_2589_final_reg_ack_1 : boolean;
  signal ptr_deref_2592_store_0_req_0 : boolean;
  signal ptr_deref_2592_store_0_ack_0 : boolean;
  signal ptr_deref_2592_store_0_req_1 : boolean;
  signal ptr_deref_2592_store_0_ack_1 : boolean;
  signal type_cast_2601_inst_req_0 : boolean;
  signal type_cast_2601_inst_ack_0 : boolean;
  signal type_cast_2601_inst_req_1 : boolean;
  signal type_cast_2601_inst_ack_1 : boolean;
  signal type_cast_2665_inst_req_0 : boolean;
  signal type_cast_2665_inst_ack_0 : boolean;
  signal type_cast_2665_inst_req_1 : boolean;
  signal type_cast_2665_inst_ack_1 : boolean;
  signal array_obj_ref_2671_index_offset_req_0 : boolean;
  signal array_obj_ref_2671_index_offset_ack_0 : boolean;
  signal array_obj_ref_2671_index_offset_req_1 : boolean;
  signal array_obj_ref_2671_index_offset_ack_1 : boolean;
  signal addr_of_2672_final_reg_req_0 : boolean;
  signal addr_of_2672_final_reg_ack_0 : boolean;
  signal addr_of_2672_final_reg_req_1 : boolean;
  signal addr_of_2672_final_reg_ack_1 : boolean;
  signal type_cast_2458_inst_req_1 : boolean;
  signal type_cast_2458_inst_ack_1 : boolean;
  signal phi_stmt_2453_req_1 : boolean;
  signal type_cast_2464_inst_req_0 : boolean;
  signal type_cast_2464_inst_ack_0 : boolean;
  signal type_cast_2464_inst_req_1 : boolean;
  signal type_cast_2464_inst_ack_1 : boolean;
  signal phi_stmt_2459_req_1 : boolean;
  signal type_cast_2449_inst_req_0 : boolean;
  signal type_cast_2449_inst_ack_0 : boolean;
  signal type_cast_2449_inst_req_1 : boolean;
  signal type_cast_2449_inst_ack_1 : boolean;
  signal phi_stmt_2446_req_0 : boolean;
  signal type_cast_2456_inst_req_0 : boolean;
  signal type_cast_2456_inst_ack_0 : boolean;
  signal type_cast_2456_inst_req_1 : boolean;
  signal type_cast_2456_inst_ack_1 : boolean;
  signal phi_stmt_2453_req_0 : boolean;
  signal type_cast_2462_inst_req_0 : boolean;
  signal type_cast_2462_inst_ack_0 : boolean;
  signal type_cast_2462_inst_req_1 : boolean;
  signal type_cast_2462_inst_ack_1 : boolean;
  signal phi_stmt_2459_req_0 : boolean;
  signal phi_stmt_2446_ack_0 : boolean;
  signal phi_stmt_2453_ack_0 : boolean;
  signal phi_stmt_2459_ack_0 : boolean;
  signal phi_stmt_2786_req_1 : boolean;
  signal type_cast_2798_inst_req_0 : boolean;
  signal type_cast_2798_inst_ack_0 : boolean;
  signal type_cast_2798_inst_req_1 : boolean;
  signal type_cast_2798_inst_ack_1 : boolean;
  signal phi_stmt_2793_req_1 : boolean;
  signal type_cast_2804_inst_req_0 : boolean;
  signal type_cast_2804_inst_ack_0 : boolean;
  signal type_cast_2804_inst_req_1 : boolean;
  signal type_cast_2804_inst_ack_1 : boolean;
  signal phi_stmt_2799_req_1 : boolean;
  signal type_cast_2789_inst_req_0 : boolean;
  signal type_cast_2789_inst_ack_0 : boolean;
  signal type_cast_2789_inst_req_1 : boolean;
  signal type_cast_2789_inst_ack_1 : boolean;
  signal phi_stmt_2786_req_0 : boolean;
  signal type_cast_2796_inst_req_0 : boolean;
  signal type_cast_2796_inst_ack_0 : boolean;
  signal type_cast_2796_inst_req_1 : boolean;
  signal type_cast_2796_inst_ack_1 : boolean;
  signal phi_stmt_2793_req_0 : boolean;
  signal type_cast_2802_inst_req_0 : boolean;
  signal type_cast_2802_inst_ack_0 : boolean;
  signal type_cast_2802_inst_req_1 : boolean;
  signal type_cast_2802_inst_ack_1 : boolean;
  signal phi_stmt_2799_req_0 : boolean;
  signal phi_stmt_2786_ack_0 : boolean;
  signal phi_stmt_2793_ack_0 : boolean;
  signal phi_stmt_2799_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_D_CP_5934_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_D_CP_5934_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_D_CP_5934_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_D_CP_5934_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_D_CP_5934: Block -- control-path 
    signal zeropad3D_D_CP_5934_elements: BooleanArray(138 downto 0);
    -- 
  begin -- 
    zeropad3D_D_CP_5934_elements(0) <= zeropad3D_D_CP_5934_start;
    zeropad3D_D_CP_5934_symbol <= zeropad3D_D_CP_5934_elements(90);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/$entry
      -- CP-element group 0: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322__entry__
      -- CP-element group 0: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2301/branch_block_stmt_2301__entry__
      -- CP-element group 0: 	 branch_block_stmt_2301/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_6000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(0), ack => RPIPE_Block3_starting_2303_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	138 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	100 
    -- CP-element group 1: 	102 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	105 
    -- CP-element group 1: 	106 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_2301/merge_stmt_2785__exit__
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Update/cr
      -- 
    rr_6865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(1), ack => type_cast_2449_inst_req_0); -- 
    cr_6870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(1), ack => type_cast_2449_inst_req_1); -- 
    rr_6888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(1), ack => type_cast_2456_inst_req_0); -- 
    cr_6893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(1), ack => type_cast_2456_inst_req_1); -- 
    rr_6911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(1), ack => type_cast_2462_inst_req_0); -- 
    cr_6916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(1), ack => type_cast_2462_inst_req_1); -- 
    zeropad3D_D_CP_5934_elements(1) <= zeropad3D_D_CP_5934_elements(138);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_update_start_
      -- 
    ra_6001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2303_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(2)); -- 
    cr_6005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(2), ack => RPIPE_Block3_starting_2303_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2303_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Sample/rr
      -- 
    ca_6006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2303_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(3)); -- 
    rr_6014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(3), ack => RPIPE_Block3_starting_2306_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_sample_completed_
      -- 
    ra_6015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2306_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(4)); -- 
    cr_6019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(4), ack => RPIPE_Block3_starting_2306_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2306_Update/$exit
      -- 
    ca_6020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2306_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(5)); -- 
    rr_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(5), ack => RPIPE_Block3_starting_2309_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Update/$entry
      -- 
    ra_6029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2309_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(6)); -- 
    cr_6033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(6), ack => RPIPE_Block3_starting_2309_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2309_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Sample/$entry
      -- 
    ca_6034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2309_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(7)); -- 
    rr_6042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(7), ack => RPIPE_Block3_starting_2312_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_update_start_
      -- 
    ra_6043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2312_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(8)); -- 
    cr_6047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(8), ack => RPIPE_Block3_starting_2312_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2312_Update/$exit
      -- 
    ca_6048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2312_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(9)); -- 
    rr_6056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(9), ack => RPIPE_Block3_starting_2315_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_update_start_
      -- 
    ra_6057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2315_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(10)); -- 
    cr_6061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(10), ack => RPIPE_Block3_starting_2315_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2315_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Sample/$entry
      -- 
    ca_6062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2315_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(11)); -- 
    rr_6070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(11), ack => RPIPE_Block3_starting_2318_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Sample/$exit
      -- 
    ra_6071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2318_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(12)); -- 
    cr_6075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(12), ack => RPIPE_Block3_starting_2318_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2318_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Sample/rr
      -- 
    ca_6076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2318_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(13)); -- 
    rr_6084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(13), ack => RPIPE_Block3_starting_2321_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Update/cr
      -- 
    ra_6085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2321_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(14)); -- 
    cr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(14), ack => RPIPE_Block3_starting_2321_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	33 
    -- CP-element group 15: 	32 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15:  members (61) 
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/$exit
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443__entry__
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322__exit__
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2304_to_assign_stmt_2322/RPIPE_Block3_starting_2321_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Update/cr
      -- 
    ca_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2321_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(15)); -- 
    rr_6101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2326_inst_req_0); -- 
    cr_6106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2326_inst_req_1); -- 
    rr_6115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2336_inst_req_0); -- 
    cr_6120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2336_inst_req_1); -- 
    rr_6129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2346_inst_req_0); -- 
    cr_6134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2346_inst_req_1); -- 
    rr_6143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2350_inst_req_0); -- 
    cr_6148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2350_inst_req_1); -- 
    rr_6157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2354_inst_req_0); -- 
    cr_6162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2354_inst_req_1); -- 
    rr_6171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2358_inst_req_0); -- 
    cr_6176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2358_inst_req_1); -- 
    rr_6185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2367_inst_req_0); -- 
    cr_6190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2367_inst_req_1); -- 
    rr_6199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2371_inst_req_0); -- 
    cr_6204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2371_inst_req_1); -- 
    rr_6213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2401_inst_req_0); -- 
    cr_6218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(15), ack => type_cast_2401_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Sample/ra
      -- 
    ra_6102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2326_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2326_Update/ca
      -- 
    ca_6107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2326_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Sample/ra
      -- 
    ra_6116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2336_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2336_Update/ca
      -- 
    ca_6121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2336_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Sample/ra
      -- 
    ra_6130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2346_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2346_Update/ca
      -- 
    ca_6135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2346_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Sample/ra
      -- 
    ra_6144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2350_Update/ca
      -- 
    ca_6149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Sample/ra
      -- 
    ra_6158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2354_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2354_Update/ca
      -- 
    ca_6163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2354_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Sample/ra
      -- 
    ra_6172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2358_Update/ca
      -- 
    ca_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Sample/ra
      -- 
    ra_6186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2367_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2367_Update/ca
      -- 
    ca_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2367_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Sample/ra
      -- 
    ra_6200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2371_Update/ca
      -- 
    ca_6205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2371_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Sample/ra
      -- 
    ra_6214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/type_cast_2401_Update/ca
      -- 
    ca_6219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	19 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	91 
    -- CP-element group 34: 	92 
    -- CP-element group 34: 	93 
    -- CP-element group 34: 	95 
    -- CP-element group 34: 	96 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2446/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443__exit__
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2301/assign_stmt_2327_to_assign_stmt_2443/$exit
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Update/cr
      -- 
    rr_6816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(34), ack => type_cast_2458_inst_req_0); -- 
    cr_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(34), ack => type_cast_2458_inst_req_1); -- 
    rr_6839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(34), ack => type_cast_2464_inst_req_0); -- 
    cr_6844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(34), ack => type_cast_2464_inst_req_1); -- 
    zeropad3D_D_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(31) & zeropad3D_D_CP_5934_elements(33) & zeropad3D_D_CP_5934_elements(17) & zeropad3D_D_CP_5934_elements(19) & zeropad3D_D_CP_5934_elements(21) & zeropad3D_D_CP_5934_elements(23) & zeropad3D_D_CP_5934_elements(25) & zeropad3D_D_CP_5934_elements(27) & zeropad3D_D_CP_5934_elements(29);
      gj_zeropad3D_D_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	113 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Sample/ra
      -- 
    ra_6231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2469_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	113 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (13) 
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496__entry__
      -- CP-element group 36: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495__exit__
      -- CP-element group 36: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/$exit
      -- CP-element group 36: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_2301/R_orx_xcond_2497_place
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2301/if_stmt_2496_else_link/$entry
      -- 
    ca_6236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2469_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(36)); -- 
    branch_req_6244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(36), ack => if_stmt_2496_branch_req_0); -- 
    -- CP-element group 37:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	40 
    -- CP-element group 37:  members (18) 
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532__entry__
      -- CP-element group 37: 	 branch_block_stmt_2301/merge_stmt_2502__exit__
      -- CP-element group 37: 	 branch_block_stmt_2301/merge_stmt_2502_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_2301/if_stmt_2496_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_2301/if_stmt_2496_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_2301/whilex_xbody_lorx_xlhsx_xfalse64
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/$entry
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_2301/whilex_xbody_lorx_xlhsx_xfalse64_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_2301/whilex_xbody_lorx_xlhsx_xfalse64_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_2301/merge_stmt_2502_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_2301/merge_stmt_2502_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_2301/merge_stmt_2502_PhiAck/dummy
      -- 
    if_choice_transition_6249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2496_branch_ack_1, ack => zeropad3D_D_CP_5934_elements(37)); -- 
    rr_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(37), ack => type_cast_2506_inst_req_0); -- 
    cr_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(37), ack => type_cast_2506_inst_req_1); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	114 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_2301/if_stmt_2496_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_2301/if_stmt_2496_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_2301/whilex_xbody_ifx_xthen
      -- CP-element group 38: 	 branch_block_stmt_2301/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2301/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_6253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2496_branch_ack_0, ack => zeropad3D_D_CP_5934_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Sample/ra
      -- 
    ra_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(39)); -- 
    -- CP-element group 40:  branch  transition  place  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (13) 
      -- CP-element group 40: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532__exit__
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533__entry__
      -- CP-element group 40: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/$exit
      -- CP-element group 40: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2301/assign_stmt_2507_to_assign_stmt_2532/type_cast_2506_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533_dead_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533_eval_test/$entry
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533_eval_test/$exit
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533_eval_test/branch_req
      -- CP-element group 40: 	 branch_block_stmt_2301/R_orx_xcond194_2534_place
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533_if_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_2301/if_stmt_2533_else_link/$entry
      -- 
    ca_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(40)); -- 
    branch_req_6280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(40), ack => if_stmt_2533_branch_req_0); -- 
    -- CP-element group 41:  fork  transition  place  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	64 
    -- CP-element group 41: 	62 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	58 
    -- CP-element group 41: 	60 
    -- CP-element group 41: 	66 
    -- CP-element group 41: 	68 
    -- CP-element group 41: 	70 
    -- CP-element group 41: 	72 
    -- CP-element group 41: 	75 
    -- CP-element group 41:  members (46) 
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_complete/req
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702__entry__
      -- CP-element group 41: 	 branch_block_stmt_2301/merge_stmt_2597__exit__
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2301/merge_stmt_2597_PhiReqMerge
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_2301/if_stmt_2533_if_link/$exit
      -- CP-element group 41: 	 branch_block_stmt_2301/if_stmt_2533_if_link/if_choice_transition
      -- CP-element group 41: 	 branch_block_stmt_2301/lorx_xlhsx_xfalse64_ifx_xelse
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_complete/req
      -- CP-element group 41: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2301/lorx_xlhsx_xfalse64_ifx_xelse_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/lorx_xlhsx_xfalse64_ifx_xelse_PhiReq/$exit
      -- CP-element group 41: 	 branch_block_stmt_2301/merge_stmt_2597_PhiAck/$entry
      -- CP-element group 41: 	 branch_block_stmt_2301/merge_stmt_2597_PhiAck/$exit
      -- CP-element group 41: 	 branch_block_stmt_2301/merge_stmt_2597_PhiAck/dummy
      -- 
    if_choice_transition_6285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2533_branch_ack_1, ack => zeropad3D_D_CP_5934_elements(41)); -- 
    req_6618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => addr_of_2697_final_reg_req_1); -- 
    cr_6572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => type_cast_2690_inst_req_1); -- 
    cr_6668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => ptr_deref_2700_store_0_req_1); -- 
    req_6603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => array_obj_ref_2696_index_offset_req_1); -- 
    cr_6553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => ptr_deref_2676_load_0_req_1); -- 
    rr_6443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => type_cast_2601_inst_req_0); -- 
    cr_6448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => type_cast_2601_inst_req_1); -- 
    cr_6462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => type_cast_2665_inst_req_1); -- 
    req_6493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => array_obj_ref_2671_index_offset_req_1); -- 
    req_6508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(41), ack => addr_of_2672_final_reg_req_1); -- 
    -- CP-element group 42:  transition  place  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	114 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_2301/if_stmt_2533_else_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_2301/if_stmt_2533_else_link/else_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_2301/lorx_xlhsx_xfalse64_ifx_xthen
      -- CP-element group 42: 	 branch_block_stmt_2301/lorx_xlhsx_xfalse64_ifx_xthen_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_2301/lorx_xlhsx_xfalse64_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_6289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2533_branch_ack_0, ack => zeropad3D_D_CP_5934_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	114 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Sample/ra
      -- 
    ra_6303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2543_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	114 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Update/ca
      -- 
    ca_6308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2543_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	114 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Sample/ra
      -- 
    ra_6317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2548_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	114 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Update/ca
      -- 
    ca_6322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2548_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Sample/rr
      -- 
    rr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(47), ack => type_cast_2582_inst_req_0); -- 
    zeropad3D_D_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(44) & zeropad3D_D_CP_5934_elements(46);
      gj_zeropad3D_D_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Sample/ra
      -- 
    ra_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	114 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Sample/req
      -- 
    ca_6336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(49)); -- 
    req_6361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(49), ack => array_obj_ref_2588_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	56 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Sample/ack
      -- 
    ack_6362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2588_index_offset_ack_0, ack => zeropad3D_D_CP_5934_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	114 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_request/req
      -- 
    ack_6367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2588_index_offset_ack_1, ack => zeropad3D_D_CP_5934_elements(51)); -- 
    req_6376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(51), ack => addr_of_2589_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_request/ack
      -- 
    ack_6377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2589_final_reg_ack_0, ack => zeropad3D_D_CP_5934_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	114 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (28) 
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/ptr_deref_2592_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/ptr_deref_2592_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/ptr_deref_2592_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/ptr_deref_2592_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/word_access_start/word_0/rr
      -- 
    ack_6382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2589_final_reg_ack_1, ack => zeropad3D_D_CP_5934_elements(53)); -- 
    rr_6420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(53), ack => ptr_deref_2592_store_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Sample/word_access_start/word_0/ra
      -- 
    ra_6421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2592_store_0_ack_0, ack => zeropad3D_D_CP_5934_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	114 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/word_access_complete/word_0/ca
      -- 
    ca_6432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2592_store_0_ack_1, ack => zeropad3D_D_CP_5934_elements(55)); -- 
    -- CP-element group 56:  join  transition  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	50 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	115 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2301/ifx_xthen_ifx_xend
      -- CP-element group 56: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595__exit__
      -- CP-element group 56: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/$exit
      -- CP-element group 56: 	 branch_block_stmt_2301/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2301/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(55) & zeropad3D_D_CP_5934_elements(50);
      gj_zeropad3D_D_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Sample/ra
      -- 
    ra_6444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2601_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	67 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2601_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Sample/rr
      -- 
    ca_6449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2601_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(58)); -- 
    rr_6457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(58), ack => type_cast_2665_inst_req_0); -- 
    rr_6567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(58), ack => type_cast_2690_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Sample/ra
      -- 
    ra_6458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2665_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	41 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (16) 
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2665_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_scale_1/scale_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Sample/req
      -- 
    ca_6463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2665_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(60)); -- 
    req_6488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(60), ack => array_obj_ref_2671_index_offset_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	76 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Sample/ack
      -- 
    ack_6489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_index_offset_ack_0, ack => zeropad3D_D_CP_5934_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	41 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (11) 
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_offset_calculated
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_final_index_sum_regn_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2671_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_request/$entry
      -- CP-element group 62: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_request/req
      -- 
    ack_6494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2671_index_offset_ack_1, ack => zeropad3D_D_CP_5934_elements(62)); -- 
    req_6503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(62), ack => addr_of_2672_final_reg_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_request/$exit
      -- CP-element group 63: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_request/ack
      -- 
    ack_6504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2672_final_reg_ack_0, ack => zeropad3D_D_CP_5934_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	41 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (24) 
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_word_addrgen/$exit
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_addr_resize/base_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_word_addrgen/$entry
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/word_access_start/word_0/rr
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_addr_resize/base_resize_req
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_word_addrgen/root_register_ack
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_word_addrgen/root_register_req
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2672_complete/ack
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_word_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_address_resized
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_addr_resize/$entry
      -- CP-element group 64: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_base_addr_resize/$exit
      -- 
    ack_6509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2672_final_reg_ack_1, ack => zeropad3D_D_CP_5934_elements(64)); -- 
    rr_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(64), ack => ptr_deref_2676_load_0_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/word_access_start/word_0/ra
      -- CP-element group 65: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_sample_completed_
      -- 
    ra_6543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2676_load_0_ack_0, ack => zeropad3D_D_CP_5934_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	41 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	73 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/ptr_deref_2676_Merge/merge_ack
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/ptr_deref_2676_Merge/merge_req
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/ptr_deref_2676_Merge/$exit
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/ptr_deref_2676_Merge/$entry
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/word_access_complete/word_0/ca
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2676_update_completed_
      -- 
    ca_6554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2676_load_0_ack_1, ack => zeropad3D_D_CP_5934_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	58 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_sample_completed_
      -- 
    ra_6568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	41 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_resize_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_resize_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_computed_1
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_resize_1/index_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_scaled_1
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_scale_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_resized_1
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/type_cast_2690_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_resize_1/index_resize_req
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Sample/req
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_scale_1/scale_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_scale_1/scale_rename_req
      -- CP-element group 68: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_index_scale_1/$exit
      -- 
    ca_6573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(68)); -- 
    req_6598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(68), ack => array_obj_ref_2696_index_offset_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	76 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_sample_complete
      -- 
    ack_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2696_index_offset_ack_0, ack => zeropad3D_D_CP_5934_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	41 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (11) 
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_offset_calculated
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_request/req
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_request/$entry
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/array_obj_ref_2696_final_index_sum_regn_Update/$exit
      -- 
    ack_6604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2696_index_offset_ack_1, ack => zeropad3D_D_CP_5934_elements(70)); -- 
    req_6613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(70), ack => addr_of_2697_final_reg_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_request/ack
      -- CP-element group 71: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_request/$exit
      -- 
    ack_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2697_final_reg_ack_0, ack => zeropad3D_D_CP_5934_elements(71)); -- 
    -- CP-element group 72:  fork  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	41 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (19) 
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_word_addrgen/root_register_ack
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_complete/ack
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/addr_of_2697_complete/$exit
      -- 
    ack_6619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2697_final_reg_ack_1, ack => zeropad3D_D_CP_5934_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/ptr_deref_2700_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/ptr_deref_2700_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/ptr_deref_2700_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/ptr_deref_2700_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/word_access_start/word_0/rr
      -- 
    rr_6657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(73), ack => ptr_deref_2700_store_0_req_0); -- 
    zeropad3D_D_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(66) & zeropad3D_D_CP_5934_elements(72);
      gj_zeropad3D_D_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Sample/word_access_start/word_0/ra
      -- 
    ra_6658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2700_store_0_ack_0, ack => zeropad3D_D_CP_5934_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/word_access_complete/word_0/ca
      -- CP-element group 75: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/ptr_deref_2700_Update/$exit
      -- 
    ca_6669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2700_store_0_ack_1, ack => zeropad3D_D_CP_5934_elements(75)); -- 
    -- CP-element group 76:  join  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	61 
    -- CP-element group 76: 	69 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	115 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_2301/ifx_xelse_ifx_xend
      -- CP-element group 76: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702__exit__
      -- CP-element group 76: 	 branch_block_stmt_2301/assign_stmt_2602_to_assign_stmt_2702/$exit
      -- CP-element group 76: 	 branch_block_stmt_2301/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2301/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(61) & zeropad3D_D_CP_5934_elements(69) & zeropad3D_D_CP_5934_elements(75);
      gj_zeropad3D_D_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	115 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Sample/$exit
      -- 
    ra_6681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2708_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(77)); -- 
    -- CP-element group 78:  branch  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	115 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (13) 
      -- CP-element group 78: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723_eval_test/$entry
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723__entry__
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723_dead_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722__exit__
      -- CP-element group 78: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/$exit
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723_else_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723_if_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723_eval_test/branch_req
      -- CP-element group 78: 	 branch_block_stmt_2301/if_stmt_2723_eval_test/$exit
      -- CP-element group 78: 	 branch_block_stmt_2301/R_cmp148_2724_place
      -- 
    ca_6686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2708_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(78)); -- 
    branch_req_6694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(78), ack => if_stmt_2723_branch_req_0); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	124 
    -- CP-element group 79: 	125 
    -- CP-element group 79: 	127 
    -- CP-element group 79: 	128 
    -- CP-element group 79: 	130 
    -- CP-element group 79: 	131 
    -- CP-element group 79:  members (40) 
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188
      -- CP-element group 79: 	 branch_block_stmt_2301/assign_stmt_2735__exit__
      -- CP-element group 79: 	 branch_block_stmt_2301/assign_stmt_2735__entry__
      -- CP-element group 79: 	 branch_block_stmt_2301/merge_stmt_2729_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_2301/merge_stmt_2729__exit__
      -- CP-element group 79: 	 branch_block_stmt_2301/assign_stmt_2735/$exit
      -- CP-element group 79: 	 branch_block_stmt_2301/assign_stmt_2735/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/if_stmt_2723_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_2301/if_stmt_2723_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xend_ifx_xthen150
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xend_ifx_xthen150_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xend_ifx_xthen150_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_2301/merge_stmt_2729_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/merge_stmt_2729_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_2301/merge_stmt_2729_PhiAck/dummy
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2723_branch_ack_1, ack => zeropad3D_D_CP_5934_elements(79)); -- 
    rr_7071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(79), ack => type_cast_2789_inst_req_0); -- 
    cr_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(79), ack => type_cast_2789_inst_req_1); -- 
    rr_7094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(79), ack => type_cast_2796_inst_req_0); -- 
    cr_7099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(79), ack => type_cast_2796_inst_req_1); -- 
    rr_7117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(79), ack => type_cast_2802_inst_req_0); -- 
    cr_7122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(79), ack => type_cast_2802_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  place  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80: 	84 
    -- CP-element group 80: 	86 
    -- CP-element group 80:  members (24) 
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2301/merge_stmt_2737_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778__entry__
      -- CP-element group 80: 	 branch_block_stmt_2301/merge_stmt_2737__exit__
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_2301/if_stmt_2723_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_2301/if_stmt_2723_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_2301/ifx_xend_ifx_xelse155
      -- CP-element group 80: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/ifx_xend_ifx_xelse155_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/ifx_xend_ifx_xelse155_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_2301/merge_stmt_2737_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_2301/merge_stmt_2737_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_2301/merge_stmt_2737_PhiAck/dummy
      -- 
    else_choice_transition_6703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2723_branch_ack_0, ack => zeropad3D_D_CP_5934_elements(80)); -- 
    rr_6719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(80), ack => type_cast_2747_inst_req_0); -- 
    cr_6738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(80), ack => type_cast_2756_inst_req_1); -- 
    cr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(80), ack => type_cast_2747_inst_req_1); -- 
    cr_6752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(80), ack => type_cast_2772_inst_req_1); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_sample_completed_
      -- 
    ra_6720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2747_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2747_Update/ca
      -- 
    ca_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2747_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(82)); -- 
    rr_6733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(82), ack => type_cast_2756_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Sample/ra
      -- 
    ra_6734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2756_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Sample/$entry
      -- 
    ca_6739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(84)); -- 
    rr_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(84), ack => type_cast_2772_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Sample/$exit
      -- 
    ra_6748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(85)); -- 
    -- CP-element group 86:  branch  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	80 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (13) 
      -- CP-element group 86: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779__entry__
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/$exit
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779_else_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778__exit__
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_2301/if_stmt_2779_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2301/R_cmp180_2780_place
      -- CP-element group 86: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2301/assign_stmt_2743_to_assign_stmt_2778/type_cast_2772_Update/$exit
      -- 
    ca_6753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2772_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(86)); -- 
    branch_req_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(86), ack => if_stmt_2779_branch_req_0); -- 
    -- CP-element group 87:  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (15) 
      -- CP-element group 87: 	 branch_block_stmt_2301/assign_stmt_2812__entry__
      -- CP-element group 87: 	 branch_block_stmt_2301/merge_stmt_2807__exit__
      -- CP-element group 87: 	 branch_block_stmt_2301/merge_stmt_2807_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_2301/if_stmt_2779_if_link/if_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_2301/if_stmt_2779_if_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2301/assign_stmt_2812/$entry
      -- CP-element group 87: 	 branch_block_stmt_2301/ifx_xelse155_whilex_xend
      -- CP-element group 87: 	 branch_block_stmt_2301/ifx_xelse155_whilex_xend_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_2301/ifx_xelse155_whilex_xend_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_2301/merge_stmt_2807_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_2301/merge_stmt_2807_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_2301/merge_stmt_2807_PhiAck/dummy
      -- 
    if_choice_transition_6766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2779_branch_ack_1, ack => zeropad3D_D_CP_5934_elements(87)); -- 
    req_6783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(87), ack => WPIPE_Block3_complete_2809_inst_req_0); -- 
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	116 
    -- CP-element group 88: 	117 
    -- CP-element group 88: 	118 
    -- CP-element group 88: 	120 
    -- CP-element group 88: 	121 
    -- CP-element group 88:  members (22) 
      -- CP-element group 88: 	 branch_block_stmt_2301/if_stmt_2779_else_link/else_choice_transition
      -- CP-element group 88: 	 branch_block_stmt_2301/if_stmt_2779_else_link/$exit
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2786/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2779_branch_ack_0, ack => zeropad3D_D_CP_5934_elements(88)); -- 
    rr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(88), ack => type_cast_2798_inst_req_0); -- 
    cr_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(88), ack => type_cast_2798_inst_req_1); -- 
    rr_7045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(88), ack => type_cast_2804_inst_req_0); -- 
    cr_7050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(88), ack => type_cast_2804_inst_req_1); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Update/req
      -- CP-element group 89: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_sample_completed_
      -- 
    ack_6784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_complete_2809_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(89)); -- 
    req_6788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(89), ack => WPIPE_Block3_complete_2809_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (16) 
      -- CP-element group 90: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2301/merge_stmt_2814__exit__
      -- CP-element group 90: 	 branch_block_stmt_2301/return__
      -- CP-element group 90: 	 branch_block_stmt_2301/assign_stmt_2812__exit__
      -- CP-element group 90: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_2301/branch_block_stmt_2301__exit__
      -- CP-element group 90: 	 branch_block_stmt_2301/$exit
      -- CP-element group 90: 	 $exit
      -- CP-element group 90: 	 branch_block_stmt_2301/assign_stmt_2812/WPIPE_Block3_complete_2809_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_2301/merge_stmt_2814_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_2301/assign_stmt_2812/$exit
      -- CP-element group 90: 	 branch_block_stmt_2301/return___PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_2301/return___PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2301/merge_stmt_2814_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_2301/merge_stmt_2814_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_2301/merge_stmt_2814_PhiAck/dummy
      -- 
    ack_6789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_complete_2809_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(90)); -- 
    -- CP-element group 91:  transition  output  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	34 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_req
      -- CP-element group 91: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2452_konst_delay_trans
      -- CP-element group 91: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2446/$exit
      -- 
    phi_stmt_2446_req_6800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2446_req_6800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(91), ack => phi_stmt_2446_req_1); -- 
    -- Element group zeropad3D_D_CP_5934_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => zeropad3D_D_CP_5934_elements(34), ack => zeropad3D_D_CP_5934_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	34 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Sample/ra
      -- 
    ra_6817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2458_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	34 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/Update/ca
      -- 
    ca_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2458_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/$exit
      -- CP-element group 94: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2458/$exit
      -- CP-element group 94: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_req
      -- 
    phi_stmt_2453_req_6823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2453_req_6823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(94), ack => phi_stmt_2453_req_1); -- 
    zeropad3D_D_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(92) & zeropad3D_D_CP_5934_elements(93);
      gj_zeropad3D_D_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	34 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Sample/ra
      -- 
    ra_6840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2464_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	34 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/Update/ca
      -- 
    ca_6845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2464_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/$exit
      -- CP-element group 97: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/$exit
      -- CP-element group 97: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2464/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_req
      -- 
    phi_stmt_2459_req_6846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2459_req_6846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(97), ack => phi_stmt_2459_req_1); -- 
    zeropad3D_D_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(95) & zeropad3D_D_CP_5934_elements(96);
      gj_zeropad3D_D_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	109 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2301/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(91) & zeropad3D_D_CP_5934_elements(94) & zeropad3D_D_CP_5934_elements(97);
      gj_zeropad3D_D_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Sample/ra
      -- 
    ra_6866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2449_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/Update/ca
      -- 
    ca_6871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2449_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/$exit
      -- CP-element group 101: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/$exit
      -- CP-element group 101: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_sources/type_cast_2449/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2446/phi_stmt_2446_req
      -- 
    phi_stmt_2446_req_6872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2446_req_6872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(101), ack => phi_stmt_2446_req_0); -- 
    zeropad3D_D_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(99) & zeropad3D_D_CP_5934_elements(100);
      gj_zeropad3D_D_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Sample/ra
      -- 
    ra_6889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2456_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/Update/ca
      -- 
    ca_6894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2456_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/$exit
      -- CP-element group 104: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/$exit
      -- CP-element group 104: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_sources/type_cast_2456/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2453/phi_stmt_2453_req
      -- 
    phi_stmt_2453_req_6895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2453_req_6895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(104), ack => phi_stmt_2453_req_0); -- 
    zeropad3D_D_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(102) & zeropad3D_D_CP_5934_elements(103);
      gj_zeropad3D_D_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	1 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Sample/ra
      -- 
    ra_6912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2462_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/Update/ca
      -- 
    ca_6917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2462_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/$exit
      -- CP-element group 107: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/$exit
      -- CP-element group 107: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_sources/type_cast_2462/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/phi_stmt_2459/phi_stmt_2459_req
      -- 
    phi_stmt_2459_req_6918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2459_req_6918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(107), ack => phi_stmt_2459_req_0); -- 
    zeropad3D_D_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(105) & zeropad3D_D_CP_5934_elements(106);
      gj_zeropad3D_D_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2301/ifx_xend188_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(101) & zeropad3D_D_CP_5934_elements(104) & zeropad3D_D_CP_5934_elements(107);
      gj_zeropad3D_D_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	98 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2301/merge_stmt_2445_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_2301/merge_stmt_2445_PhiAck/$entry
      -- 
    zeropad3D_D_CP_5934_elements(109) <= OrReduce(zeropad3D_D_CP_5934_elements(98) & zeropad3D_D_CP_5934_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_2301/merge_stmt_2445_PhiAck/phi_stmt_2446_ack
      -- 
    phi_stmt_2446_ack_6923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2446_ack_0, ack => zeropad3D_D_CP_5934_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2301/merge_stmt_2445_PhiAck/phi_stmt_2453_ack
      -- 
    phi_stmt_2453_ack_6924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2453_ack_0, ack => zeropad3D_D_CP_5934_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2301/merge_stmt_2445_PhiAck/phi_stmt_2459_ack
      -- 
    phi_stmt_2459_ack_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2459_ack_0, ack => zeropad3D_D_CP_5934_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	35 
    -- CP-element group 113: 	36 
    -- CP-element group 113:  members (10) 
      -- CP-element group 113: 	 branch_block_stmt_2301/merge_stmt_2445__exit__
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495__entry__
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/$entry
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_update_start_
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_2301/assign_stmt_2470_to_assign_stmt_2495/type_cast_2469_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_2301/merge_stmt_2445_PhiAck/$exit
      -- 
    rr_6230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(113), ack => type_cast_2469_inst_req_0); -- 
    cr_6235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(113), ack => type_cast_2469_inst_req_1); -- 
    zeropad3D_D_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(110) & zeropad3D_D_CP_5934_elements(111) & zeropad3D_D_CP_5934_elements(112);
      gj_zeropad3D_D_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  merge  fork  transition  place  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	38 
    -- CP-element group 114: 	42 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	43 
    -- CP-element group 114: 	51 
    -- CP-element group 114: 	44 
    -- CP-element group 114: 	53 
    -- CP-element group 114: 	45 
    -- CP-element group 114: 	46 
    -- CP-element group 114: 	55 
    -- CP-element group 114: 	49 
    -- CP-element group 114:  members (33) 
      -- CP-element group 114: 	 branch_block_stmt_2301/merge_stmt_2539__exit__
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595__entry__
      -- CP-element group 114: 	 branch_block_stmt_2301/merge_stmt_2539_PhiReqMerge
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2543_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2548_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/type_cast_2582_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_update_start
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/array_obj_ref_2588_final_index_sum_regn_Update/req
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/addr_of_2589_complete/req
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/word_access_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/word_access_complete/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/assign_stmt_2544_to_assign_stmt_2595/ptr_deref_2592_Update/word_access_complete/word_0/cr
      -- CP-element group 114: 	 branch_block_stmt_2301/merge_stmt_2539_PhiAck/$entry
      -- CP-element group 114: 	 branch_block_stmt_2301/merge_stmt_2539_PhiAck/$exit
      -- CP-element group 114: 	 branch_block_stmt_2301/merge_stmt_2539_PhiAck/dummy
      -- 
    rr_6302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => type_cast_2543_inst_req_0); -- 
    cr_6307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => type_cast_2543_inst_req_1); -- 
    rr_6316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => type_cast_2548_inst_req_0); -- 
    cr_6321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => type_cast_2548_inst_req_1); -- 
    cr_6335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => type_cast_2582_inst_req_1); -- 
    req_6366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => array_obj_ref_2588_index_offset_req_1); -- 
    req_6381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => addr_of_2589_final_reg_req_1); -- 
    cr_6431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(114), ack => ptr_deref_2592_store_0_req_1); -- 
    zeropad3D_D_CP_5934_elements(114) <= OrReduce(zeropad3D_D_CP_5934_elements(38) & zeropad3D_D_CP_5934_elements(42));
    -- CP-element group 115:  merge  fork  transition  place  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	56 
    -- CP-element group 115: 	76 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	77 
    -- CP-element group 115: 	78 
    -- CP-element group 115:  members (13) 
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_2301/merge_stmt_2704_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_update_start_
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722__entry__
      -- CP-element group 115: 	 branch_block_stmt_2301/merge_stmt_2704__exit__
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/type_cast_2708_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_2301/assign_stmt_2709_to_assign_stmt_2722/$entry
      -- CP-element group 115: 	 branch_block_stmt_2301/merge_stmt_2704_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_2301/merge_stmt_2704_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_2301/merge_stmt_2704_PhiAck/dummy
      -- 
    cr_6685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(115), ack => type_cast_2708_inst_req_1); -- 
    rr_6680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(115), ack => type_cast_2708_inst_req_0); -- 
    zeropad3D_D_CP_5934_elements(115) <= OrReduce(zeropad3D_D_CP_5934_elements(56) & zeropad3D_D_CP_5934_elements(76));
    -- CP-element group 116:  transition  output  delay-element  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	88 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	123 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2786/$exit
      -- CP-element group 116: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2792_konst_delay_trans
      -- CP-element group 116: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_req
      -- 
    phi_stmt_2786_req_7006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2786_req_7006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(116), ack => phi_stmt_2786_req_1); -- 
    -- Element group zeropad3D_D_CP_5934_elements(116) is a control-delay.
    cp_element_116_delay: control_delay_element  generic map(name => " 116_delay", delay_value => 1)  port map(req => zeropad3D_D_CP_5934_elements(88), ack => zeropad3D_D_CP_5934_elements(116), clk => clk, reset =>reset);
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	88 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Sample/ra
      -- 
    ra_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2798_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/Update/ca
      -- 
    ca_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2798_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/$exit
      -- CP-element group 119: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/$exit
      -- CP-element group 119: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2798/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_req
      -- 
    phi_stmt_2793_req_7029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2793_req_7029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(119), ack => phi_stmt_2793_req_1); -- 
    zeropad3D_D_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(117) & zeropad3D_D_CP_5934_elements(118);
      gj_zeropad3D_D_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	88 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Sample/ra
      -- 
    ra_7046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2804_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	88 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/Update/ca
      -- 
    ca_7051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2804_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/$exit
      -- CP-element group 122: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/$exit
      -- CP-element group 122: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2804/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_req
      -- 
    phi_stmt_2799_req_7052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2799_req_7052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(122), ack => phi_stmt_2799_req_1); -- 
    zeropad3D_D_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(120) & zeropad3D_D_CP_5934_elements(121);
      gj_zeropad3D_D_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	116 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	134 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2301/ifx_xelse155_ifx_xend188_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(116) & zeropad3D_D_CP_5934_elements(119) & zeropad3D_D_CP_5934_elements(122);
      gj_zeropad3D_D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	79 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Sample/ra
      -- 
    ra_7072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2789_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/Update/ca
      -- 
    ca_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2789_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	133 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/$exit
      -- CP-element group 126: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/$exit
      -- CP-element group 126: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_sources/type_cast_2789/SplitProtocol/$exit
      -- CP-element group 126: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2786/phi_stmt_2786_req
      -- 
    phi_stmt_2786_req_7078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2786_req_7078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(126), ack => phi_stmt_2786_req_0); -- 
    zeropad3D_D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(124) & zeropad3D_D_CP_5934_elements(125);
      gj_zeropad3D_D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	79 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Sample/ra
      -- 
    ra_7095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2796_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	79 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/Update/ca
      -- 
    ca_7100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2796_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/$exit
      -- CP-element group 129: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/$exit
      -- CP-element group 129: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/$exit
      -- CP-element group 129: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_sources/type_cast_2796/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2793/phi_stmt_2793_req
      -- 
    phi_stmt_2793_req_7101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2793_req_7101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(129), ack => phi_stmt_2793_req_0); -- 
    zeropad3D_D_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(127) & zeropad3D_D_CP_5934_elements(128);
      gj_zeropad3D_D_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	79 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Sample/ra
      -- 
    ra_7118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_0, ack => zeropad3D_D_CP_5934_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	79 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/Update/ca
      -- 
    ca_7123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2802_inst_ack_1, ack => zeropad3D_D_CP_5934_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/$exit
      -- CP-element group 132: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/$exit
      -- CP-element group 132: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/$exit
      -- CP-element group 132: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_sources/type_cast_2802/SplitProtocol/$exit
      -- CP-element group 132: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/phi_stmt_2799/phi_stmt_2799_req
      -- 
    phi_stmt_2799_req_7124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2799_req_7124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5934_elements(132), ack => phi_stmt_2799_req_0); -- 
    zeropad3D_D_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(130) & zeropad3D_D_CP_5934_elements(131);
      gj_zeropad3D_D_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	126 
    -- CP-element group 133: 	129 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_2301/ifx_xthen150_ifx_xend188_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(126) & zeropad3D_D_CP_5934_elements(129) & zeropad3D_D_CP_5934_elements(132);
      gj_zeropad3D_D_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  merge  fork  transition  place  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	123 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2301/merge_stmt_2785_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_2301/merge_stmt_2785_PhiAck/$entry
      -- 
    zeropad3D_D_CP_5934_elements(134) <= OrReduce(zeropad3D_D_CP_5934_elements(123) & zeropad3D_D_CP_5934_elements(133));
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_2301/merge_stmt_2785_PhiAck/phi_stmt_2786_ack
      -- 
    phi_stmt_2786_ack_7129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2786_ack_0, ack => zeropad3D_D_CP_5934_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_2301/merge_stmt_2785_PhiAck/phi_stmt_2793_ack
      -- 
    phi_stmt_2793_ack_7130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2793_ack_0, ack => zeropad3D_D_CP_5934_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_2301/merge_stmt_2785_PhiAck/phi_stmt_2799_ack
      -- 
    phi_stmt_2799_ack_7131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2799_ack_0, ack => zeropad3D_D_CP_5934_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	1 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_2301/merge_stmt_2785_PhiAck/$exit
      -- 
    zeropad3D_D_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5934_elements(135) & zeropad3D_D_CP_5934_elements(136) & zeropad3D_D_CP_5934_elements(137);
      gj_zeropad3D_D_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5934_elements(138), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2385_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2441_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2576_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2659_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2684_wire : std_logic_vector(31 downto 0);
    signal R_idxprom135_2670_resized : std_logic_vector(13 downto 0);
    signal R_idxprom135_2670_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom140_2695_resized : std_logic_vector(13 downto 0);
    signal R_idxprom140_2695_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2587_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2587_scaled : std_logic_vector(13 downto 0);
    signal add107_2627 : std_logic_vector(31 downto 0);
    signal add116_2632 : std_logic_vector(31 downto 0);
    signal add126_2647 : std_logic_vector(31 downto 0);
    signal add132_2652 : std_logic_vector(31 downto 0);
    signal add145_2715 : std_logic_vector(31 downto 0);
    signal add153_2735 : std_logic_vector(15 downto 0);
    signal add163_2398 : std_logic_vector(31 downto 0);
    signal add179_2413 : std_logic_vector(31 downto 0);
    signal add78_2423 : std_logic_vector(31 downto 0);
    signal add89_2564 : std_logic_vector(31 downto 0);
    signal add95_2569 : std_logic_vector(31 downto 0);
    signal add_2418 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2588_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2588_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2588_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2588_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2588_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2588_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2671_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2671_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2671_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2671_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2671_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2671_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2696_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2696_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2696_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2696_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2696_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2696_root_address : std_logic_vector(13 downto 0);
    signal arrayidx136_2673 : std_logic_vector(31 downto 0);
    signal arrayidx141_2698 : std_logic_vector(31 downto 0);
    signal arrayidx_2590 : std_logic_vector(31 downto 0);
    signal call1_2307 : std_logic_vector(7 downto 0);
    signal call2_2310 : std_logic_vector(7 downto 0);
    signal call3_2313 : std_logic_vector(7 downto 0);
    signal call4_2316 : std_logic_vector(7 downto 0);
    signal call5_2319 : std_logic_vector(7 downto 0);
    signal call6_2322 : std_logic_vector(7 downto 0);
    signal call_2304 : std_logic_vector(7 downto 0);
    signal cmp148_2722 : std_logic_vector(0 downto 0);
    signal cmp164_2753 : std_logic_vector(0 downto 0);
    signal cmp180_2778 : std_logic_vector(0 downto 0);
    signal cmp62_2490 : std_logic_vector(0 downto 0);
    signal cmp69_2514 : std_logic_vector(0 downto 0);
    signal cmp69x_xnot_2520 : std_logic_vector(0 downto 0);
    signal cmp79_2527 : std_logic_vector(0 downto 0);
    signal cmp_2477 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_2483 : std_logic_vector(0 downto 0);
    signal conv109_2443 : std_logic_vector(31 downto 0);
    signal conv10_2337 : std_logic_vector(15 downto 0);
    signal conv144_2709 : std_logic_vector(31 downto 0);
    signal conv158_2748 : std_logic_vector(31 downto 0);
    signal conv172_2773 : std_logic_vector(31 downto 0);
    signal conv174_2402 : std_logic_vector(31 downto 0);
    signal conv36_2347 : std_logic_vector(31 downto 0);
    signal conv38_2351 : std_logic_vector(31 downto 0);
    signal conv42_2355 : std_logic_vector(31 downto 0);
    signal conv44_2359 : std_logic_vector(31 downto 0);
    signal conv51_2470 : std_logic_vector(31 downto 0);
    signal conv53_2368 : std_logic_vector(31 downto 0);
    signal conv66_2507 : std_logic_vector(31 downto 0);
    signal conv83_2544 : std_logic_vector(31 downto 0);
    signal conv85_2372 : std_logic_vector(31 downto 0);
    signal conv87_2549 : std_logic_vector(31 downto 0);
    signal conv91_2387 : std_logic_vector(31 downto 0);
    signal conv99_2602 : std_logic_vector(31 downto 0);
    signal conv_2327 : std_logic_vector(15 downto 0);
    signal div11_2343 : std_logic_vector(15 downto 0);
    signal div175_2408 : std_logic_vector(31 downto 0);
    signal div_2333 : std_logic_vector(15 downto 0);
    signal idxprom135_2666 : std_logic_vector(63 downto 0);
    signal idxprom140_2691 : std_logic_vector(63 downto 0);
    signal idxprom_2583 : std_logic_vector(63 downto 0);
    signal inc169_2757 : std_logic_vector(15 downto 0);
    signal inc169x_xix_x2_2762 : std_logic_vector(15 downto 0);
    signal inc_2743 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_2793 : std_logic_vector(15 downto 0);
    signal ix_x2_2453 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_2799 : std_logic_vector(15 downto 0);
    signal jx_x1_2459 : std_logic_vector(15 downto 0);
    signal jx_x2_2768 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_2786 : std_logic_vector(15 downto 0);
    signal kx_x1_2446 : std_logic_vector(15 downto 0);
    signal mul106_2612 : std_logic_vector(31 downto 0);
    signal mul115_2622 : std_logic_vector(31 downto 0);
    signal mul125_2637 : std_logic_vector(31 downto 0);
    signal mul131_2642 : std_logic_vector(31 downto 0);
    signal mul45_2364 : std_logic_vector(31 downto 0);
    signal mul88_2554 : std_logic_vector(31 downto 0);
    signal mul94_2559 : std_logic_vector(31 downto 0);
    signal mul_2429 : std_logic_vector(31 downto 0);
    signal orx_xcond194_2532 : std_logic_vector(0 downto 0);
    signal orx_xcond_2495 : std_logic_vector(0 downto 0);
    signal ptr_deref_2592_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2592_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2592_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2592_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2592_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2592_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2676_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2676_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2676_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2676_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2676_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2700_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2700_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2700_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2700_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2700_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2700_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext193_2378 : std_logic_vector(31 downto 0);
    signal sext_2434 : std_logic_vector(31 downto 0);
    signal shl_2393 : std_logic_vector(31 downto 0);
    signal shr134_2661 : std_logic_vector(31 downto 0);
    signal shr139_2686 : std_logic_vector(31 downto 0);
    signal shr_2578 : std_logic_vector(31 downto 0);
    signal sub114_2617 : std_logic_vector(31 downto 0);
    signal sub_2607 : std_logic_vector(31 downto 0);
    signal tmp137_2677 : std_logic_vector(63 downto 0);
    signal type_cast_2331_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2341_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2376_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2381_wire : std_logic_vector(31 downto 0);
    signal type_cast_2384_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2391_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2406_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2427_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2437_wire : std_logic_vector(31 downto 0);
    signal type_cast_2440_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2449_wire : std_logic_vector(15 downto 0);
    signal type_cast_2452_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2456_wire : std_logic_vector(15 downto 0);
    signal type_cast_2458_wire : std_logic_vector(15 downto 0);
    signal type_cast_2462_wire : std_logic_vector(15 downto 0);
    signal type_cast_2464_wire : std_logic_vector(15 downto 0);
    signal type_cast_2468_wire : std_logic_vector(31 downto 0);
    signal type_cast_2473_wire : std_logic_vector(31 downto 0);
    signal type_cast_2475_wire : std_logic_vector(31 downto 0);
    signal type_cast_2481_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2486_wire : std_logic_vector(31 downto 0);
    signal type_cast_2488_wire : std_logic_vector(31 downto 0);
    signal type_cast_2505_wire : std_logic_vector(31 downto 0);
    signal type_cast_2510_wire : std_logic_vector(31 downto 0);
    signal type_cast_2512_wire : std_logic_vector(31 downto 0);
    signal type_cast_2518_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2523_wire : std_logic_vector(31 downto 0);
    signal type_cast_2525_wire : std_logic_vector(31 downto 0);
    signal type_cast_2542_wire : std_logic_vector(31 downto 0);
    signal type_cast_2547_wire : std_logic_vector(31 downto 0);
    signal type_cast_2572_wire : std_logic_vector(31 downto 0);
    signal type_cast_2575_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2581_wire : std_logic_vector(63 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2600_wire : std_logic_vector(31 downto 0);
    signal type_cast_2655_wire : std_logic_vector(31 downto 0);
    signal type_cast_2658_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2664_wire : std_logic_vector(63 downto 0);
    signal type_cast_2680_wire : std_logic_vector(31 downto 0);
    signal type_cast_2683_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2689_wire : std_logic_vector(63 downto 0);
    signal type_cast_2707_wire : std_logic_vector(31 downto 0);
    signal type_cast_2713_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2718_wire : std_logic_vector(31 downto 0);
    signal type_cast_2720_wire : std_logic_vector(31 downto 0);
    signal type_cast_2733_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2741_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2746_wire : std_logic_vector(31 downto 0);
    signal type_cast_2771_wire : std_logic_vector(31 downto 0);
    signal type_cast_2789_wire : std_logic_vector(15 downto 0);
    signal type_cast_2792_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2796_wire : std_logic_vector(15 downto 0);
    signal type_cast_2798_wire : std_logic_vector(15 downto 0);
    signal type_cast_2802_wire : std_logic_vector(15 downto 0);
    signal type_cast_2804_wire : std_logic_vector(15 downto 0);
    signal type_cast_2811_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_2588_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2588_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2588_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2588_resized_base_address <= "00000000000000";
    array_obj_ref_2671_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2671_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2671_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2671_resized_base_address <= "00000000000000";
    array_obj_ref_2696_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2696_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2696_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2696_resized_base_address <= "00000000000000";
    ptr_deref_2592_word_offset_0 <= "00000000000000";
    ptr_deref_2676_word_offset_0 <= "00000000000000";
    ptr_deref_2700_word_offset_0 <= "00000000000000";
    type_cast_2331_wire_constant <= "0000000000000001";
    type_cast_2341_wire_constant <= "0000000000000010";
    type_cast_2376_wire_constant <= "00000000000000000000000000010000";
    type_cast_2384_wire_constant <= "00000000000000000000000000010000";
    type_cast_2391_wire_constant <= "00000000000000000000000000000001";
    type_cast_2406_wire_constant <= "00000000000000000000000000000001";
    type_cast_2427_wire_constant <= "00000000000000000000000000010000";
    type_cast_2440_wire_constant <= "00000000000000000000000000010000";
    type_cast_2452_wire_constant <= "0000000000000000";
    type_cast_2481_wire_constant <= "1";
    type_cast_2518_wire_constant <= "1";
    type_cast_2575_wire_constant <= "00000000000000000000000000000010";
    type_cast_2594_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2658_wire_constant <= "00000000000000000000000000000010";
    type_cast_2683_wire_constant <= "00000000000000000000000000000010";
    type_cast_2713_wire_constant <= "00000000000000000000000000000100";
    type_cast_2733_wire_constant <= "0000000000000100";
    type_cast_2741_wire_constant <= "0000000000000001";
    type_cast_2792_wire_constant <= "0000000000000000";
    type_cast_2811_wire_constant <= "00000001";
    phi_stmt_2446: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2449_wire & type_cast_2452_wire_constant;
      req <= phi_stmt_2446_req_0 & phi_stmt_2446_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2446",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2446_ack_0,
          idata => idata,
          odata => kx_x1_2446,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2446
    phi_stmt_2453: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2456_wire & type_cast_2458_wire;
      req <= phi_stmt_2453_req_0 & phi_stmt_2453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2453",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2453_ack_0,
          idata => idata,
          odata => ix_x2_2453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2453
    phi_stmt_2459: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2462_wire & type_cast_2464_wire;
      req <= phi_stmt_2459_req_0 & phi_stmt_2459_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2459",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2459_ack_0,
          idata => idata,
          odata => jx_x1_2459,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2459
    phi_stmt_2786: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2789_wire & type_cast_2792_wire_constant;
      req <= phi_stmt_2786_req_0 & phi_stmt_2786_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2786",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2786_ack_0,
          idata => idata,
          odata => kx_x0x_xph_2786,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2786
    phi_stmt_2793: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2796_wire & type_cast_2798_wire;
      req <= phi_stmt_2793_req_0 & phi_stmt_2793_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2793",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2793_ack_0,
          idata => idata,
          odata => ix_x1x_xph_2793,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2793
    phi_stmt_2799: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2802_wire & type_cast_2804_wire;
      req <= phi_stmt_2799_req_0 & phi_stmt_2799_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2799",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2799_ack_0,
          idata => idata,
          odata => jx_x0x_xph_2799,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2799
    -- flow-through select operator MUX_2767_inst
    jx_x2_2768 <= div_2333 when (cmp164_2753(0) /=  '0') else inc_2743;
    addr_of_2589_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2589_final_reg_req_0;
      addr_of_2589_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2589_final_reg_req_1;
      addr_of_2589_final_reg_ack_1<= rack(0);
      addr_of_2589_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2589_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2588_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2672_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2672_final_reg_req_0;
      addr_of_2672_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2672_final_reg_req_1;
      addr_of_2672_final_reg_ack_1<= rack(0);
      addr_of_2672_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2672_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2671_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx136_2673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2697_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2697_final_reg_req_0;
      addr_of_2697_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2697_final_reg_req_1;
      addr_of_2697_final_reg_ack_1<= rack(0);
      addr_of_2697_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2697_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2696_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx141_2698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2326_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2326_inst_req_0;
      type_cast_2326_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2326_inst_req_1;
      type_cast_2326_inst_ack_1<= rack(0);
      type_cast_2326_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2326_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2327,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2336_inst_req_0;
      type_cast_2336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2336_inst_req_1;
      type_cast_2336_inst_ack_1<= rack(0);
      type_cast_2336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_2337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2346_inst_req_0;
      type_cast_2346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2346_inst_req_1;
      type_cast_2346_inst_ack_1<= rack(0);
      type_cast_2346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_2310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_2347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2350_inst_req_0;
      type_cast_2350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2350_inst_req_1;
      type_cast_2350_inst_ack_1<= rack(0);
      type_cast_2350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_2351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2354_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2354_inst_req_0;
      type_cast_2354_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2354_inst_req_1;
      type_cast_2354_inst_ack_1<= rack(0);
      type_cast_2354_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2354_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_2319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_2355,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2358_inst_req_0;
      type_cast_2358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2358_inst_req_1;
      type_cast_2358_inst_ack_1<= rack(0);
      type_cast_2358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_2316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_2359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2367_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2367_inst_req_0;
      type_cast_2367_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2367_inst_req_1;
      type_cast_2367_inst_ack_1<= rack(0);
      type_cast_2367_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2367_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_2322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_2368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2371_inst_req_0;
      type_cast_2371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2371_inst_req_1;
      type_cast_2371_inst_ack_1<= rack(0);
      type_cast_2371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_2319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2381_inst
    process(sext193_2378) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext193_2378(31 downto 0);
      type_cast_2381_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2386_inst
    process(ASHR_i32_i32_2385_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2385_wire(31 downto 0);
      conv91_2387 <= tmp_var; -- 
    end process;
    type_cast_2401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2401_inst_req_0;
      type_cast_2401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2401_inst_req_1;
      type_cast_2401_inst_ack_1<= rack(0);
      type_cast_2401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv174_2402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2437_inst
    process(sext_2434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2434(31 downto 0);
      type_cast_2437_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2442_inst
    process(ASHR_i32_i32_2441_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2441_wire(31 downto 0);
      conv109_2443 <= tmp_var; -- 
    end process;
    type_cast_2449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2449_inst_req_0;
      type_cast_2449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2449_inst_req_1;
      type_cast_2449_inst_ack_1<= rack(0);
      type_cast_2449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_2786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2449_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2456_inst_req_0;
      type_cast_2456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2456_inst_req_1;
      type_cast_2456_inst_ack_1<= rack(0);
      type_cast_2456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_2793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2456_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2458_inst_req_0;
      type_cast_2458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2458_inst_req_1;
      type_cast_2458_inst_ack_1<= rack(0);
      type_cast_2458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div11_2343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2458_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2462_inst_req_0;
      type_cast_2462_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2462_inst_req_1;
      type_cast_2462_inst_ack_1<= rack(0);
      type_cast_2462_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2462_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_2799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2462_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2464_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2464_inst_req_0;
      type_cast_2464_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2464_inst_req_1;
      type_cast_2464_inst_ack_1<= rack(0);
      type_cast_2464_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2464_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2464_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2469_inst_req_0;
      type_cast_2469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2469_inst_req_1;
      type_cast_2469_inst_ack_1<= rack(0);
      type_cast_2469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2468_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_2470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2473_inst
    process(conv51_2470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv51_2470(31 downto 0);
      type_cast_2473_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2475_inst
    process(conv53_2368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_2368(31 downto 0);
      type_cast_2475_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2486_inst
    process(conv51_2470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv51_2470(31 downto 0);
      type_cast_2486_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2488_inst
    process(add_2418) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_2418(31 downto 0);
      type_cast_2488_wire <= tmp_var; -- 
    end process;
    type_cast_2506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2506_inst_req_0;
      type_cast_2506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2506_inst_req_1;
      type_cast_2506_inst_ack_1<= rack(0);
      type_cast_2506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2505_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2507,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2510_inst
    process(conv66_2507) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv66_2507(31 downto 0);
      type_cast_2510_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2512_inst
    process(conv53_2368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_2368(31 downto 0);
      type_cast_2512_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2523_inst
    process(conv66_2507) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv66_2507(31 downto 0);
      type_cast_2523_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2525_inst
    process(add78_2423) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add78_2423(31 downto 0);
      type_cast_2525_wire <= tmp_var; -- 
    end process;
    type_cast_2543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2543_inst_req_0;
      type_cast_2543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2543_inst_req_1;
      type_cast_2543_inst_ack_1<= rack(0);
      type_cast_2543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2542_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_2544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2548_inst_req_0;
      type_cast_2548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2548_inst_req_1;
      type_cast_2548_inst_ack_1<= rack(0);
      type_cast_2548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2547_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_2549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2572_inst
    process(add95_2569) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add95_2569(31 downto 0);
      type_cast_2572_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2577_inst
    process(ASHR_i32_i32_2576_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2576_wire(31 downto 0);
      shr_2578 <= tmp_var; -- 
    end process;
    type_cast_2582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2582_inst_req_0;
      type_cast_2582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2582_inst_req_1;
      type_cast_2582_inst_ack_1<= rack(0);
      type_cast_2582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2581_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2601_inst_req_0;
      type_cast_2601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2601_inst_req_1;
      type_cast_2601_inst_ack_1<= rack(0);
      type_cast_2601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2600_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2655_inst
    process(add116_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add116_2632(31 downto 0);
      type_cast_2655_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2660_inst
    process(ASHR_i32_i32_2659_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2659_wire(31 downto 0);
      shr134_2661 <= tmp_var; -- 
    end process;
    type_cast_2665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2665_inst_req_0;
      type_cast_2665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2665_inst_req_1;
      type_cast_2665_inst_ack_1<= rack(0);
      type_cast_2665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2664_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom135_2666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2680_inst
    process(add132_2652) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add132_2652(31 downto 0);
      type_cast_2680_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2685_inst
    process(ASHR_i32_i32_2684_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2684_wire(31 downto 0);
      shr139_2686 <= tmp_var; -- 
    end process;
    type_cast_2690_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2690_inst_req_0;
      type_cast_2690_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2690_inst_req_1;
      type_cast_2690_inst_ack_1<= rack(0);
      type_cast_2690_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2690_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2689_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom140_2691,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2708_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2708_inst_req_0;
      type_cast_2708_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2708_inst_req_1;
      type_cast_2708_inst_ack_1<= rack(0);
      type_cast_2708_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2708_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2707_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_2709,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2718_inst
    process(add145_2715) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add145_2715(31 downto 0);
      type_cast_2718_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2720_inst
    process(conv36_2347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_2347(31 downto 0);
      type_cast_2720_wire <= tmp_var; -- 
    end process;
    type_cast_2747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2747_inst_req_0;
      type_cast_2747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2747_inst_req_1;
      type_cast_2747_inst_ack_1<= rack(0);
      type_cast_2747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2746_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_2748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2756_inst_req_0;
      type_cast_2756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2756_inst_req_1;
      type_cast_2756_inst_ack_1<= rack(0);
      type_cast_2756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp164_2753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc169_2757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2772_inst_req_0;
      type_cast_2772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2772_inst_req_1;
      type_cast_2772_inst_ack_1<= rack(0);
      type_cast_2772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2771_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv172_2773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2789_inst_req_0;
      type_cast_2789_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2789_inst_req_1;
      type_cast_2789_inst_ack_1<= rack(0);
      type_cast_2789_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2789_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add153_2735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2789_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2796_inst_req_0;
      type_cast_2796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2796_inst_req_1;
      type_cast_2796_inst_ack_1<= rack(0);
      type_cast_2796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_2453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2796_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2798_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2798_inst_req_0;
      type_cast_2798_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2798_inst_req_1;
      type_cast_2798_inst_ack_1<= rack(0);
      type_cast_2798_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2798_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc169x_xix_x2_2762,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2798_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2802_inst_req_0;
      type_cast_2802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2802_inst_req_1;
      type_cast_2802_inst_ack_1<= rack(0);
      type_cast_2802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_2459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2802_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2804_inst_req_0;
      type_cast_2804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2804_inst_req_1;
      type_cast_2804_inst_ack_1<= rack(0);
      type_cast_2804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_2768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2804_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2588_index_1_rename
    process(R_idxprom_2587_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2587_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2587_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2588_index_1_resize
    process(idxprom_2583) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2583;
      ov := iv(13 downto 0);
      R_idxprom_2587_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2588_root_address_inst
    process(array_obj_ref_2588_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2588_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2588_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2671_index_1_rename
    process(R_idxprom135_2670_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom135_2670_resized;
      ov(13 downto 0) := iv;
      R_idxprom135_2670_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2671_index_1_resize
    process(idxprom135_2666) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom135_2666;
      ov := iv(13 downto 0);
      R_idxprom135_2670_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2671_root_address_inst
    process(array_obj_ref_2671_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2671_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2671_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2696_index_1_rename
    process(R_idxprom140_2695_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom140_2695_resized;
      ov(13 downto 0) := iv;
      R_idxprom140_2695_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2696_index_1_resize
    process(idxprom140_2691) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom140_2691;
      ov := iv(13 downto 0);
      R_idxprom140_2695_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2696_root_address_inst
    process(array_obj_ref_2696_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2696_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2696_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2592_addr_0
    process(ptr_deref_2592_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2592_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2592_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2592_base_resize
    process(arrayidx_2590) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2590;
      ov := iv(13 downto 0);
      ptr_deref_2592_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2592_gather_scatter
    process(type_cast_2594_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2594_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2592_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2592_root_address_inst
    process(ptr_deref_2592_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2592_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2592_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2676_addr_0
    process(ptr_deref_2676_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2676_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2676_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2676_base_resize
    process(arrayidx136_2673) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx136_2673;
      ov := iv(13 downto 0);
      ptr_deref_2676_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2676_gather_scatter
    process(ptr_deref_2676_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2676_data_0;
      ov(63 downto 0) := iv;
      tmp137_2677 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2676_root_address_inst
    process(ptr_deref_2676_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2676_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2676_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2700_addr_0
    process(ptr_deref_2700_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2700_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2700_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2700_base_resize
    process(arrayidx141_2698) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx141_2698;
      ov := iv(13 downto 0);
      ptr_deref_2700_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2700_gather_scatter
    process(tmp137_2677) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp137_2677;
      ov(63 downto 0) := iv;
      ptr_deref_2700_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2700_root_address_inst
    process(ptr_deref_2700_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2700_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2700_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2496_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_2495;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2496_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2496_branch_req_0,
          ack0 => if_stmt_2496_branch_ack_0,
          ack1 => if_stmt_2496_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2533_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond194_2532;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2533_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2533_branch_req_0,
          ack0 => if_stmt_2533_branch_ack_0,
          ack1 => if_stmt_2533_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2723_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp148_2722;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2723_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2723_branch_req_0,
          ack0 => if_stmt_2723_branch_ack_0,
          ack1 => if_stmt_2723_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2779_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp180_2778;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2779_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2779_branch_req_0,
          ack0 => if_stmt_2779_branch_ack_0,
          ack1 => if_stmt_2779_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2734_inst
    process(kx_x1_2446) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_2446, type_cast_2733_wire_constant, tmp_var);
      add153_2735 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2742_inst
    process(jx_x1_2459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_2459, type_cast_2741_wire_constant, tmp_var);
      inc_2743 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2761_inst
    process(inc169_2757, ix_x2_2453) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc169_2757, ix_x2_2453, tmp_var);
      inc169x_xix_x2_2762 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2397_inst
    process(shl_2393, conv38_2351) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_2393, conv38_2351, tmp_var);
      add163_2398 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2412_inst
    process(shl_2393, div175_2408) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_2393, div175_2408, tmp_var);
      add179_2413 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2417_inst
    process(conv53_2368, div175_2408) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv53_2368, div175_2408, tmp_var);
      add_2418 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2422_inst
    process(conv53_2368, conv38_2351) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv53_2368, conv38_2351, tmp_var);
      add78_2423 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2563_inst
    process(mul94_2559, conv83_2544) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul94_2559, conv83_2544, tmp_var);
      add89_2564 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2568_inst
    process(add89_2564, mul88_2554) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add89_2564, mul88_2554, tmp_var);
      add95_2569 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2626_inst
    process(mul115_2622, conv99_2602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul115_2622, conv99_2602, tmp_var);
      add107_2627 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2631_inst
    process(add107_2627, mul106_2612) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add107_2627, mul106_2612, tmp_var);
      add116_2632 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2646_inst
    process(mul131_2642, conv99_2602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul131_2642, conv99_2602, tmp_var);
      add126_2647 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2651_inst
    process(add126_2647, mul125_2637) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add126_2647, mul125_2637, tmp_var);
      add132_2652 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2714_inst
    process(conv144_2709) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv144_2709, type_cast_2713_wire_constant, tmp_var);
      add145_2715 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2494_inst
    process(cmpx_xnot_2483, cmp62_2490) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_2483, cmp62_2490, tmp_var);
      orx_xcond_2495 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2531_inst
    process(cmp69x_xnot_2520, cmp79_2527) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp69x_xnot_2520, cmp79_2527, tmp_var);
      orx_xcond194_2532 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2385_inst
    process(type_cast_2381_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2381_wire, type_cast_2384_wire_constant, tmp_var);
      ASHR_i32_i32_2385_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2441_inst
    process(type_cast_2437_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2437_wire, type_cast_2440_wire_constant, tmp_var);
      ASHR_i32_i32_2441_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2576_inst
    process(type_cast_2572_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2572_wire, type_cast_2575_wire_constant, tmp_var);
      ASHR_i32_i32_2576_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2659_inst
    process(type_cast_2655_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2655_wire, type_cast_2658_wire_constant, tmp_var);
      ASHR_i32_i32_2659_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2684_inst
    process(type_cast_2680_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2680_wire, type_cast_2683_wire_constant, tmp_var);
      ASHR_i32_i32_2684_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2752_inst
    process(conv158_2748, add163_2398) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv158_2748, add163_2398, tmp_var);
      cmp164_2753 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2777_inst
    process(conv172_2773, add179_2413) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv172_2773, add179_2413, tmp_var);
      cmp180_2778 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2332_inst
    process(conv_2327) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_2327, type_cast_2331_wire_constant, tmp_var);
      div_2333 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2342_inst
    process(conv10_2337) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv10_2337, type_cast_2341_wire_constant, tmp_var);
      div11_2343 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2407_inst
    process(conv174_2402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv174_2402, type_cast_2406_wire_constant, tmp_var);
      div175_2408 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2363_inst
    process(conv42_2355, conv44_2359) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_2355, conv44_2359, tmp_var);
      mul45_2364 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2433_inst
    process(mul_2429, conv36_2347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_2429, conv36_2347, tmp_var);
      sext_2434 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2553_inst
    process(conv87_2549, conv85_2372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv87_2549, conv85_2372, tmp_var);
      mul88_2554 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2558_inst
    process(conv51_2470, conv91_2387) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv51_2470, conv91_2387, tmp_var);
      mul94_2559 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2611_inst
    process(sub_2607, conv36_2347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_2607, conv36_2347, tmp_var);
      mul106_2612 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2621_inst
    process(sub114_2617, conv109_2443) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub114_2617, conv109_2443, tmp_var);
      mul115_2622 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2636_inst
    process(conv66_2507, conv85_2372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv66_2507, conv85_2372, tmp_var);
      mul125_2637 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2641_inst
    process(conv51_2470, conv91_2387) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv51_2470, conv91_2387, tmp_var);
      mul131_2642 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2377_inst
    process(mul45_2364) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul45_2364, type_cast_2376_wire_constant, tmp_var);
      sext193_2378 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2392_inst
    process(conv53_2368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_2368, type_cast_2391_wire_constant, tmp_var);
      shl_2393 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2428_inst
    process(conv38_2351) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv38_2351, type_cast_2427_wire_constant, tmp_var);
      mul_2429 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2476_inst
    process(type_cast_2473_wire, type_cast_2475_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2473_wire, type_cast_2475_wire, tmp_var);
      cmp_2477 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2489_inst
    process(type_cast_2486_wire, type_cast_2488_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2486_wire, type_cast_2488_wire, tmp_var);
      cmp62_2490 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2513_inst
    process(type_cast_2510_wire, type_cast_2512_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2510_wire, type_cast_2512_wire, tmp_var);
      cmp69_2514 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2526_inst
    process(type_cast_2523_wire, type_cast_2525_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2523_wire, type_cast_2525_wire, tmp_var);
      cmp79_2527 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2721_inst
    process(type_cast_2718_wire, type_cast_2720_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2718_wire, type_cast_2720_wire, tmp_var);
      cmp148_2722 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2606_inst
    process(conv66_2507, conv53_2368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv66_2507, conv53_2368, tmp_var);
      sub_2607 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2616_inst
    process(conv51_2470, conv53_2368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv51_2470, conv53_2368, tmp_var);
      sub114_2617 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2482_inst
    process(cmp_2477) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_2477, type_cast_2481_wire_constant, tmp_var);
      cmpx_xnot_2483 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2519_inst
    process(cmp69_2514) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp69_2514, type_cast_2518_wire_constant, tmp_var);
      cmp69x_xnot_2520 <= tmp_var; --
    end process;
    -- shared split operator group (46) : array_obj_ref_2588_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2587_scaled;
      array_obj_ref_2588_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2588_index_offset_req_0;
      array_obj_ref_2588_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2588_index_offset_req_1;
      array_obj_ref_2588_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_2671_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom135_2670_scaled;
      array_obj_ref_2671_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2671_index_offset_req_0;
      array_obj_ref_2671_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2671_index_offset_req_1;
      array_obj_ref_2671_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_2696_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom140_2695_scaled;
      array_obj_ref_2696_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2696_index_offset_req_0;
      array_obj_ref_2696_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2696_index_offset_req_1;
      array_obj_ref_2696_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- unary operator type_cast_2468_inst
    process(ix_x2_2453) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_2453, tmp_var);
      type_cast_2468_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2505_inst
    process(jx_x1_2459) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2459, tmp_var);
      type_cast_2505_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2542_inst
    process(kx_x1_2446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2446, tmp_var);
      type_cast_2542_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2547_inst
    process(jx_x1_2459) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2459, tmp_var);
      type_cast_2547_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2581_inst
    process(shr_2578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2578, tmp_var);
      type_cast_2581_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2600_inst
    process(kx_x1_2446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2446, tmp_var);
      type_cast_2600_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2664_inst
    process(shr134_2661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr134_2661, tmp_var);
      type_cast_2664_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2689_inst
    process(shr139_2686) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr139_2686, tmp_var);
      type_cast_2689_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2707_inst
    process(kx_x1_2446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2446, tmp_var);
      type_cast_2707_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2746_inst
    process(inc_2743) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2743, tmp_var);
      type_cast_2746_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2771_inst
    process(inc169x_xix_x2_2762) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc169x_xix_x2_2762, tmp_var);
      type_cast_2771_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2676_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2676_load_0_req_0;
      ptr_deref_2676_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2676_load_0_req_1;
      ptr_deref_2676_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2676_word_address_0;
      ptr_deref_2676_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2592_store_0 ptr_deref_2700_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2592_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2700_store_0_req_0;
      ptr_deref_2592_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2700_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2592_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2700_store_0_req_1;
      ptr_deref_2592_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2700_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2592_word_address_0 & ptr_deref_2700_word_address_0;
      data_in <= ptr_deref_2592_data_0 & ptr_deref_2700_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_starting_2303_inst RPIPE_Block3_starting_2306_inst RPIPE_Block3_starting_2309_inst RPIPE_Block3_starting_2312_inst RPIPE_Block3_starting_2315_inst RPIPE_Block3_starting_2318_inst RPIPE_Block3_starting_2321_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block3_starting_2303_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_starting_2306_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_starting_2309_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_starting_2312_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_starting_2315_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_starting_2318_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_starting_2321_inst_req_0;
      RPIPE_Block3_starting_2303_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_starting_2306_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_starting_2309_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_starting_2312_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_starting_2315_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_starting_2318_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_starting_2321_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block3_starting_2303_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_starting_2306_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_starting_2309_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_starting_2312_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_starting_2315_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_starting_2318_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_starting_2321_inst_req_1;
      RPIPE_Block3_starting_2303_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_starting_2306_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_starting_2309_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_starting_2312_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_starting_2315_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_starting_2318_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_starting_2321_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call_2304 <= data_out(55 downto 48);
      call1_2307 <= data_out(47 downto 40);
      call2_2310 <= data_out(39 downto 32);
      call3_2313 <= data_out(31 downto 24);
      call4_2316 <= data_out(23 downto 16);
      call5_2319 <= data_out(15 downto 8);
      call6_2322 <= data_out(7 downto 0);
      Block3_starting_read_0_gI: SplitGuardInterface generic map(name => "Block3_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block3_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_starting_pipe_read_req(0),
          oack => Block3_starting_pipe_read_ack(0),
          odata => Block3_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_complete_2809_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_complete_2809_inst_req_0;
      WPIPE_Block3_complete_2809_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_complete_2809_inst_req_1;
      WPIPE_Block3_complete_2809_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2811_wire_constant;
      Block3_complete_write_0_gI: SplitGuardInterface generic map(name => "Block3_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_complete_pipe_write_req(0),
          oack => Block3_complete_pipe_write_ack(0),
          odata => Block3_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_E is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block4_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block4_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block4_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block4_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block4_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block4_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_E;
architecture zeropad3D_E_arch of zeropad3D_E is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_E_CP_7148_start: Boolean;
  signal zeropad3D_E_CP_7148_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block4_starting_2829_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2835_inst_ack_0 : boolean;
  signal type_cast_2865_inst_req_1 : boolean;
  signal type_cast_2861_inst_req_0 : boolean;
  signal type_cast_2874_inst_req_1 : boolean;
  signal type_cast_2874_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2835_inst_req_1 : boolean;
  signal type_cast_2874_inst_req_0 : boolean;
  signal type_cast_2874_inst_ack_0 : boolean;
  signal type_cast_2843_inst_ack_0 : boolean;
  signal type_cast_2865_inst_ack_1 : boolean;
  signal type_cast_2865_inst_req_0 : boolean;
  signal type_cast_2865_inst_ack_0 : boolean;
  signal type_cast_2861_inst_req_1 : boolean;
  signal type_cast_2861_inst_ack_1 : boolean;
  signal type_cast_2853_inst_req_0 : boolean;
  signal RPIPE_Block4_starting_2832_inst_req_1 : boolean;
  signal RPIPE_Block4_starting_2832_inst_ack_1 : boolean;
  signal type_cast_2853_inst_ack_0 : boolean;
  signal type_cast_2843_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2838_inst_req_0 : boolean;
  signal RPIPE_Block4_starting_2835_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2826_inst_req_0 : boolean;
  signal RPIPE_Block4_starting_2826_inst_ack_0 : boolean;
  signal type_cast_2843_inst_req_1 : boolean;
  signal RPIPE_Block4_starting_2838_inst_ack_1 : boolean;
  signal type_cast_2857_inst_req_0 : boolean;
  signal type_cast_2857_inst_req_1 : boolean;
  signal RPIPE_Block4_starting_2820_inst_req_0 : boolean;
  signal type_cast_2853_inst_req_1 : boolean;
  signal type_cast_2853_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2820_inst_ack_0 : boolean;
  signal type_cast_2857_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2838_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2826_inst_ack_1 : boolean;
  signal type_cast_2861_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2838_inst_req_1 : boolean;
  signal type_cast_2857_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2829_inst_req_0 : boolean;
  signal RPIPE_Block4_starting_2823_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2832_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2823_inst_req_1 : boolean;
  signal type_cast_2914_inst_req_1 : boolean;
  signal type_cast_2914_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2832_inst_req_0 : boolean;
  signal type_cast_3063_inst_req_0 : boolean;
  signal type_cast_3063_inst_ack_0 : boolean;
  signal type_cast_3063_inst_req_1 : boolean;
  signal type_cast_3063_inst_ack_1 : boolean;
  signal type_cast_3068_inst_req_0 : boolean;
  signal type_cast_3068_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2835_inst_req_0 : boolean;
  signal type_cast_2878_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2823_inst_ack_0 : boolean;
  signal RPIPE_Block4_starting_2823_inst_req_0 : boolean;
  signal type_cast_3026_inst_req_0 : boolean;
  signal type_cast_3026_inst_ack_0 : boolean;
  signal type_cast_3026_inst_req_1 : boolean;
  signal RPIPE_Block4_starting_2826_inst_req_1 : boolean;
  signal if_stmt_3016_branch_ack_0 : boolean;
  signal if_stmt_3053_branch_ack_1 : boolean;
  signal if_stmt_3053_branch_ack_0 : boolean;
  signal type_cast_2989_inst_req_1 : boolean;
  signal if_stmt_3016_branch_ack_1 : boolean;
  signal type_cast_3026_inst_ack_1 : boolean;
  signal if_stmt_3053_branch_req_0 : boolean;
  signal type_cast_2878_inst_req_1 : boolean;
  signal RPIPE_Block4_starting_2829_inst_ack_1 : boolean;
  signal type_cast_2989_inst_req_0 : boolean;
  signal type_cast_2989_inst_ack_0 : boolean;
  signal type_cast_2989_inst_ack_1 : boolean;
  signal RPIPE_Block4_starting_2829_inst_req_1 : boolean;
  signal type_cast_2914_inst_ack_0 : boolean;
  signal type_cast_2914_inst_req_0 : boolean;
  signal RPIPE_Block4_starting_2820_inst_ack_1 : boolean;
  signal type_cast_2843_inst_req_0 : boolean;
  signal type_cast_2878_inst_req_0 : boolean;
  signal type_cast_2878_inst_ack_0 : boolean;
  signal if_stmt_3016_branch_req_0 : boolean;
  signal RPIPE_Block4_starting_2820_inst_req_1 : boolean;
  signal type_cast_3068_inst_req_1 : boolean;
  signal type_cast_3068_inst_ack_1 : boolean;
  signal type_cast_3102_inst_req_0 : boolean;
  signal type_cast_3102_inst_ack_0 : boolean;
  signal type_cast_3102_inst_req_1 : boolean;
  signal type_cast_3102_inst_ack_1 : boolean;
  signal array_obj_ref_3108_index_offset_req_0 : boolean;
  signal array_obj_ref_3108_index_offset_ack_0 : boolean;
  signal array_obj_ref_3108_index_offset_req_1 : boolean;
  signal array_obj_ref_3108_index_offset_ack_1 : boolean;
  signal addr_of_3109_final_reg_req_0 : boolean;
  signal addr_of_3109_final_reg_ack_0 : boolean;
  signal addr_of_3109_final_reg_req_1 : boolean;
  signal addr_of_3109_final_reg_ack_1 : boolean;
  signal ptr_deref_3112_store_0_req_0 : boolean;
  signal ptr_deref_3112_store_0_ack_0 : boolean;
  signal ptr_deref_3112_store_0_req_1 : boolean;
  signal ptr_deref_3112_store_0_ack_1 : boolean;
  signal type_cast_3121_inst_req_0 : boolean;
  signal type_cast_3121_inst_ack_0 : boolean;
  signal type_cast_3121_inst_req_1 : boolean;
  signal type_cast_3121_inst_ack_1 : boolean;
  signal type_cast_3185_inst_req_0 : boolean;
  signal type_cast_3185_inst_ack_0 : boolean;
  signal type_cast_3185_inst_req_1 : boolean;
  signal type_cast_3185_inst_ack_1 : boolean;
  signal array_obj_ref_3191_index_offset_req_0 : boolean;
  signal array_obj_ref_3191_index_offset_ack_0 : boolean;
  signal array_obj_ref_3191_index_offset_req_1 : boolean;
  signal array_obj_ref_3191_index_offset_ack_1 : boolean;
  signal addr_of_3192_final_reg_req_0 : boolean;
  signal addr_of_3192_final_reg_ack_0 : boolean;
  signal addr_of_3192_final_reg_req_1 : boolean;
  signal addr_of_3192_final_reg_ack_1 : boolean;
  signal ptr_deref_3196_load_0_req_0 : boolean;
  signal ptr_deref_3196_load_0_ack_0 : boolean;
  signal ptr_deref_3196_load_0_req_1 : boolean;
  signal ptr_deref_3196_load_0_ack_1 : boolean;
  signal type_cast_3210_inst_req_0 : boolean;
  signal type_cast_3210_inst_ack_0 : boolean;
  signal type_cast_3210_inst_req_1 : boolean;
  signal type_cast_3210_inst_ack_1 : boolean;
  signal array_obj_ref_3216_index_offset_req_0 : boolean;
  signal array_obj_ref_3216_index_offset_ack_0 : boolean;
  signal array_obj_ref_3216_index_offset_req_1 : boolean;
  signal array_obj_ref_3216_index_offset_ack_1 : boolean;
  signal addr_of_3217_final_reg_req_0 : boolean;
  signal addr_of_3217_final_reg_ack_0 : boolean;
  signal addr_of_3217_final_reg_req_1 : boolean;
  signal addr_of_3217_final_reg_ack_1 : boolean;
  signal ptr_deref_3220_store_0_req_0 : boolean;
  signal ptr_deref_3220_store_0_ack_0 : boolean;
  signal ptr_deref_3220_store_0_req_1 : boolean;
  signal ptr_deref_3220_store_0_ack_1 : boolean;
  signal type_cast_3228_inst_req_0 : boolean;
  signal type_cast_3228_inst_ack_0 : boolean;
  signal type_cast_3228_inst_req_1 : boolean;
  signal type_cast_3228_inst_ack_1 : boolean;
  signal if_stmt_3243_branch_req_0 : boolean;
  signal if_stmt_3243_branch_ack_1 : boolean;
  signal if_stmt_3243_branch_ack_0 : boolean;
  signal type_cast_3267_inst_req_0 : boolean;
  signal type_cast_3267_inst_ack_0 : boolean;
  signal type_cast_3267_inst_req_1 : boolean;
  signal type_cast_3267_inst_ack_1 : boolean;
  signal type_cast_3276_inst_req_0 : boolean;
  signal type_cast_3276_inst_ack_0 : boolean;
  signal type_cast_3276_inst_req_1 : boolean;
  signal type_cast_3276_inst_ack_1 : boolean;
  signal type_cast_3293_inst_req_0 : boolean;
  signal type_cast_3293_inst_ack_0 : boolean;
  signal type_cast_3293_inst_req_1 : boolean;
  signal type_cast_3293_inst_ack_1 : boolean;
  signal if_stmt_3300_branch_req_0 : boolean;
  signal if_stmt_3300_branch_ack_1 : boolean;
  signal if_stmt_3300_branch_ack_0 : boolean;
  signal WPIPE_Block4_complete_3330_inst_req_0 : boolean;
  signal WPIPE_Block4_complete_3330_inst_ack_0 : boolean;
  signal WPIPE_Block4_complete_3330_inst_req_1 : boolean;
  signal WPIPE_Block4_complete_3330_inst_ack_1 : boolean;
  signal phi_stmt_2965_req_0 : boolean;
  signal type_cast_2975_inst_req_0 : boolean;
  signal type_cast_2975_inst_ack_0 : boolean;
  signal type_cast_2975_inst_req_1 : boolean;
  signal type_cast_2975_inst_ack_1 : boolean;
  signal phi_stmt_2972_req_0 : boolean;
  signal phi_stmt_2978_req_0 : boolean;
  signal type_cast_2971_inst_req_0 : boolean;
  signal type_cast_2971_inst_ack_0 : boolean;
  signal type_cast_2971_inst_req_1 : boolean;
  signal type_cast_2971_inst_ack_1 : boolean;
  signal phi_stmt_2965_req_1 : boolean;
  signal type_cast_2977_inst_req_0 : boolean;
  signal type_cast_2977_inst_ack_0 : boolean;
  signal type_cast_2977_inst_req_1 : boolean;
  signal type_cast_2977_inst_ack_1 : boolean;
  signal phi_stmt_2972_req_1 : boolean;
  signal type_cast_2984_inst_req_0 : boolean;
  signal type_cast_2984_inst_ack_0 : boolean;
  signal type_cast_2984_inst_req_1 : boolean;
  signal type_cast_2984_inst_ack_1 : boolean;
  signal phi_stmt_2978_req_1 : boolean;
  signal phi_stmt_2965_ack_0 : boolean;
  signal phi_stmt_2972_ack_0 : boolean;
  signal phi_stmt_2978_ack_0 : boolean;
  signal type_cast_3325_inst_req_0 : boolean;
  signal type_cast_3325_inst_ack_0 : boolean;
  signal type_cast_3325_inst_req_1 : boolean;
  signal type_cast_3325_inst_ack_1 : boolean;
  signal phi_stmt_3320_req_1 : boolean;
  signal type_cast_3319_inst_req_0 : boolean;
  signal type_cast_3319_inst_ack_0 : boolean;
  signal type_cast_3319_inst_req_1 : boolean;
  signal type_cast_3319_inst_ack_1 : boolean;
  signal phi_stmt_3314_req_1 : boolean;
  signal phi_stmt_3307_req_1 : boolean;
  signal type_cast_3323_inst_req_0 : boolean;
  signal type_cast_3323_inst_ack_0 : boolean;
  signal type_cast_3323_inst_req_1 : boolean;
  signal type_cast_3323_inst_ack_1 : boolean;
  signal phi_stmt_3320_req_0 : boolean;
  signal type_cast_3317_inst_req_0 : boolean;
  signal type_cast_3317_inst_ack_0 : boolean;
  signal type_cast_3317_inst_req_1 : boolean;
  signal type_cast_3317_inst_ack_1 : boolean;
  signal phi_stmt_3314_req_0 : boolean;
  signal type_cast_3310_inst_req_0 : boolean;
  signal type_cast_3310_inst_ack_0 : boolean;
  signal type_cast_3310_inst_req_1 : boolean;
  signal type_cast_3310_inst_ack_1 : boolean;
  signal phi_stmt_3307_req_0 : boolean;
  signal phi_stmt_3307_ack_0 : boolean;
  signal phi_stmt_3314_ack_0 : boolean;
  signal phi_stmt_3320_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_E_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_E_CP_7148_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_E_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_E_CP_7148_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_E_CP_7148_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_E_CP_7148_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_E_CP_7148: Block -- control-path 
    signal zeropad3D_E_CP_7148_elements: BooleanArray(134 downto 0);
    -- 
  begin -- 
    zeropad3D_E_CP_7148_elements(0) <= zeropad3D_E_CP_7148_start;
    zeropad3D_E_CP_7148_symbol <= zeropad3D_E_CP_7148_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2818/$entry
      -- CP-element group 0: 	 branch_block_stmt_2818/branch_block_stmt_2818__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839__entry__
      -- CP-element group 0: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/$entry
      -- 
    rr_7214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(0), ack => RPIPE_Block4_starting_2820_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	134 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	102 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2818/merge_stmt_3306__exit__
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Update/cr
      -- 
    rr_8050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(1), ack => type_cast_2971_inst_req_0); -- 
    cr_8055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(1), ack => type_cast_2971_inst_req_1); -- 
    rr_8073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(1), ack => type_cast_2977_inst_req_0); -- 
    cr_8078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(1), ack => type_cast_2977_inst_req_1); -- 
    rr_8096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(1), ack => type_cast_2984_inst_req_0); -- 
    cr_8101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(1), ack => type_cast_2984_inst_req_1); -- 
    zeropad3D_E_CP_7148_elements(1) <= zeropad3D_E_CP_7148_elements(134);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Update/cr
      -- 
    ra_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2820_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(2)); -- 
    cr_7219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(2), ack => RPIPE_Block4_starting_2820_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2820_Update/ca
      -- 
    ca_7220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2820_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(3)); -- 
    rr_7228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(3), ack => RPIPE_Block4_starting_2823_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_sample_completed_
      -- 
    ra_7229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2823_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(4)); -- 
    cr_7233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(4), ack => RPIPE_Block4_starting_2823_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2823_update_completed_
      -- 
    ca_7234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2823_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(5)); -- 
    rr_7242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(5), ack => RPIPE_Block4_starting_2826_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Update/cr
      -- 
    ra_7243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2826_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(6)); -- 
    cr_7247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(6), ack => RPIPE_Block4_starting_2826_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2826_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Sample/$entry
      -- 
    ca_7248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2826_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(7)); -- 
    rr_7256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(7), ack => RPIPE_Block4_starting_2829_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_update_start_
      -- 
    ra_7257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2829_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(8)); -- 
    cr_7261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(8), ack => RPIPE_Block4_starting_2829_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2829_Update/$exit
      -- 
    ca_7262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2829_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(9)); -- 
    rr_7270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(9), ack => RPIPE_Block4_starting_2832_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_sample_completed_
      -- 
    ra_7271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2832_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(10)); -- 
    cr_7275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(10), ack => RPIPE_Block4_starting_2832_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2832_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Sample/$entry
      -- 
    ca_7276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2832_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(11)); -- 
    rr_7284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(11), ack => RPIPE_Block4_starting_2835_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Sample/$exit
      -- 
    ra_7285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2835_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(12)); -- 
    cr_7289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(12), ack => RPIPE_Block4_starting_2835_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2835_update_completed_
      -- 
    ca_7290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2835_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(13)); -- 
    rr_7298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(13), ack => RPIPE_Block4_starting_2838_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_update_start_
      -- 
    ra_7299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2838_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(14)); -- 
    cr_7303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(14), ack => RPIPE_Block4_starting_2838_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15:  members (55) 
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962__entry__
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839__exit__
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/$exit
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2821_to_assign_stmt_2839/RPIPE_Block4_starting_2838_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Update/$entry
      -- 
    ca_7304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block4_starting_2838_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(15)); -- 
    cr_7376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2865_inst_req_1); -- 
    rr_7357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2861_inst_req_0); -- 
    cr_7390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2874_inst_req_1); -- 
    rr_7385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2874_inst_req_0); -- 
    rr_7371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2865_inst_req_0); -- 
    cr_7362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2861_inst_req_1); -- 
    rr_7329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2853_inst_req_0); -- 
    cr_7320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2843_inst_req_1); -- 
    rr_7343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2857_inst_req_0); -- 
    cr_7348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2857_inst_req_1); -- 
    cr_7334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2853_inst_req_1); -- 
    cr_7418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2914_inst_req_1); -- 
    cr_7404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2878_inst_req_1); -- 
    rr_7413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2914_inst_req_0); -- 
    rr_7315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2843_inst_req_0); -- 
    rr_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(15), ack => type_cast_2878_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Sample/$exit
      -- 
    ra_7316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2843_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2843_Update/$exit
      -- 
    ca_7321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2843_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Sample/$exit
      -- 
    ra_7330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2853_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2853_Update/ca
      -- 
    ca_7335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2853_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Sample/ra
      -- 
    ra_7344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2857_Update/ca
      -- 
    ca_7349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Sample/$exit
      -- 
    ra_7358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2861_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2861_update_completed_
      -- 
    ca_7363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2861_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_sample_completed_
      -- 
    ra_7372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2865_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2865_Update/ca
      -- 
    ca_7377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2865_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_sample_completed_
      -- 
    ra_7386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2874_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2874_Update/$exit
      -- 
    ca_7391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2874_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Sample/ra
      -- 
    ra_7400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2878_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2878_Update/$exit
      -- 
    ca_7405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2878_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Sample/$exit
      -- 
    ra_7414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/type_cast_2914_update_completed_
      -- 
    ca_7419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	21 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	25 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: 	90 
    -- CP-element group 32: 	91 
    -- CP-element group 32: 	93 
    -- CP-element group 32:  members (16) 
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody
      -- CP-element group 32: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962__exit__
      -- CP-element group 32: 	 branch_block_stmt_2818/assign_stmt_2844_to_assign_stmt_2962/$exit
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2965/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2978/$entry
      -- CP-element group 32: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/$entry
      -- 
    rr_8016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(32), ack => type_cast_2975_inst_req_0); -- 
    cr_8021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(32), ack => type_cast_2975_inst_req_1); -- 
    zeropad3D_E_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(17) & zeropad3D_E_CP_7148_elements(19) & zeropad3D_E_CP_7148_elements(21) & zeropad3D_E_CP_7148_elements(23) & zeropad3D_E_CP_7148_elements(25) & zeropad3D_E_CP_7148_elements(27) & zeropad3D_E_CP_7148_elements(29) & zeropad3D_E_CP_7148_elements(31);
      gj_zeropad3D_E_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	109 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Sample/ra
      -- 
    ra_7431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2989_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	109 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (13) 
      -- CP-element group 34: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015__exit__
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016__entry__
      -- CP-element group 34: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/$exit
      -- CP-element group 34: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016_else_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_2818/R_orx_xcond_3017_place
      -- CP-element group 34: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_2818/if_stmt_3016_eval_test/branch_req
      -- 
    ca_7436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2989_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(34)); -- 
    branch_req_7444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(34), ack => if_stmt_3016_branch_req_0); -- 
    -- CP-element group 35:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (18) 
      -- CP-element group 35: 	 branch_block_stmt_2818/merge_stmt_3022__exit__
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052__entry__
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_2818/whilex_xbody_lorx_xlhsx_xfalse60
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/$entry
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_update_start_
      -- CP-element group 35: 	 branch_block_stmt_2818/if_stmt_3016_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_2818/if_stmt_3016_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_2818/whilex_xbody_lorx_xlhsx_xfalse60_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_2818/whilex_xbody_lorx_xlhsx_xfalse60_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_2818/merge_stmt_3022_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_2818/merge_stmt_3022_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_2818/merge_stmt_3022_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_2818/merge_stmt_3022_PhiAck/dummy
      -- 
    if_choice_transition_7449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3016_branch_ack_1, ack => zeropad3D_E_CP_7148_elements(35)); -- 
    rr_7466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(35), ack => type_cast_3026_inst_req_0); -- 
    cr_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(35), ack => type_cast_3026_inst_req_1); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	110 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_2818/whilex_xbody_ifx_xthen
      -- CP-element group 36: 	 branch_block_stmt_2818/if_stmt_3016_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_2818/if_stmt_3016_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_2818/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_2818/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_7453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3016_branch_ack_0, ack => zeropad3D_E_CP_7148_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_sample_completed_
      -- 
    ra_7467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3026_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (13) 
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053__entry__
      -- CP-element group 38: 	 branch_block_stmt_2818/R_orx_xcond193_3054_place
      -- CP-element group 38: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052__exit__
      -- CP-element group 38: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053_if_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053_else_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/$exit
      -- CP-element group 38: 	 branch_block_stmt_2818/assign_stmt_3027_to_assign_stmt_3052/type_cast_3026_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_2818/if_stmt_3053_eval_test/branch_req
      -- 
    ca_7472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3026_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(38)); -- 
    branch_req_7480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(38), ack => if_stmt_3053_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222__entry__
      -- CP-element group 39: 	 branch_block_stmt_2818/lorx_xlhsx_xfalse60_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_2818/merge_stmt_3117__exit__
      -- CP-element group 39: 	 branch_block_stmt_2818/if_stmt_3053_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_2818/if_stmt_3053_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_complete/req
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_complete/req
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_update_start_
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_2818/lorx_xlhsx_xfalse60_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/lorx_xlhsx_xfalse60_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_2818/merge_stmt_3117_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_2818/merge_stmt_3117_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_2818/merge_stmt_3117_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_2818/merge_stmt_3117_PhiAck/dummy
      -- 
    if_choice_transition_7485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3053_branch_ack_1, ack => zeropad3D_E_CP_7148_elements(39)); -- 
    rr_7643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => type_cast_3121_inst_req_0); -- 
    cr_7648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => type_cast_3121_inst_req_1); -- 
    cr_7662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => type_cast_3185_inst_req_1); -- 
    req_7693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => array_obj_ref_3191_index_offset_req_1); -- 
    req_7708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => addr_of_3192_final_reg_req_1); -- 
    cr_7753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => ptr_deref_3196_load_0_req_1); -- 
    cr_7772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => type_cast_3210_inst_req_1); -- 
    req_7803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => array_obj_ref_3216_index_offset_req_1); -- 
    req_7818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => addr_of_3217_final_reg_req_1); -- 
    cr_7868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(39), ack => ptr_deref_3220_store_0_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	110 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_2818/lorx_xlhsx_xfalse60_ifx_xthen
      -- CP-element group 40: 	 branch_block_stmt_2818/if_stmt_3053_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_2818/if_stmt_3053_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_2818/lorx_xlhsx_xfalse60_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_2818/lorx_xlhsx_xfalse60_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_7489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3053_branch_ack_0, ack => zeropad3D_E_CP_7148_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	110 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_sample_completed_
      -- 
    ra_7503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3063_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	110 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Update/ca
      -- 
    ca_7508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3063_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	110 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Sample/ra
      -- 
    ra_7517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3068_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Update/ca
      -- 
    ca_7522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3068_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Sample/rr
      -- 
    rr_7530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(45), ack => type_cast_3102_inst_req_0); -- 
    zeropad3D_E_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(42) & zeropad3D_E_CP_7148_elements(44);
      gj_zeropad3D_E_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Sample/ra
      -- 
    ra_7531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3102_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	110 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_computed_1
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Sample/req
      -- 
    ca_7536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3102_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(47)); -- 
    req_7561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(47), ack => array_obj_ref_3108_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Sample/ack
      -- 
    ack_7562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3108_index_offset_ack_0, ack => zeropad3D_E_CP_7148_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	110 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_request/req
      -- 
    ack_7567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3108_index_offset_ack_1, ack => zeropad3D_E_CP_7148_elements(49)); -- 
    req_7576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(49), ack => addr_of_3109_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_request/$exit
      -- CP-element group 50: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_request/ack
      -- 
    ack_7577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3109_final_reg_ack_0, ack => zeropad3D_E_CP_7148_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	110 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_word_addrgen/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/ptr_deref_3112_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/ptr_deref_3112_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/ptr_deref_3112_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/ptr_deref_3112_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/word_access_start/word_0/rr
      -- 
    ack_7582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3109_final_reg_ack_1, ack => zeropad3D_E_CP_7148_elements(51)); -- 
    rr_7620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(51), ack => ptr_deref_3112_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Sample/word_access_start/word_0/ra
      -- 
    ra_7621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3112_store_0_ack_0, ack => zeropad3D_E_CP_7148_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	110 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/word_access_complete/word_0/ca
      -- 
    ca_7632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3112_store_0_ack_1, ack => zeropad3D_E_CP_7148_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: 	48 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	111 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2818/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115__exit__
      -- CP-element group 54: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/$exit
      -- CP-element group 54: 	 branch_block_stmt_2818/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2818/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_E_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(53) & zeropad3D_E_CP_7148_elements(48);
      gj_zeropad3D_E_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Sample/ra
      -- 
    ra_7644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3121_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3121_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Sample/rr
      -- 
    ca_7649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3121_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(56)); -- 
    rr_7657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(56), ack => type_cast_3185_inst_req_0); -- 
    rr_7767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(56), ack => type_cast_3210_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Sample/ra
      -- 
    ra_7658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3185_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3185_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Sample/req
      -- 
    ca_7663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3185_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(58)); -- 
    req_7688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(58), ack => array_obj_ref_3191_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Sample/ack
      -- 
    ack_7689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3191_index_offset_ack_0, ack => zeropad3D_E_CP_7148_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3191_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_request/req
      -- 
    ack_7694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3191_index_offset_ack_1, ack => zeropad3D_E_CP_7148_elements(60)); -- 
    req_7703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(60), ack => addr_of_3192_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_request/ack
      -- 
    ack_7704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3192_final_reg_ack_0, ack => zeropad3D_E_CP_7148_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3192_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/word_access_start/word_0/rr
      -- 
    ack_7709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3192_final_reg_ack_1, ack => zeropad3D_E_CP_7148_elements(62)); -- 
    rr_7742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(62), ack => ptr_deref_3196_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Sample/word_access_start/word_0/ra
      -- 
    ra_7743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3196_load_0_ack_0, ack => zeropad3D_E_CP_7148_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/ptr_deref_3196_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/ptr_deref_3196_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/ptr_deref_3196_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3196_Update/ptr_deref_3196_Merge/merge_ack
      -- 
    ca_7754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3196_load_0_ack_1, ack => zeropad3D_E_CP_7148_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Sample/ra
      -- 
    ra_7768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3210_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/type_cast_3210_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_computed_1
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Sample/req
      -- 
    ca_7773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3210_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(66)); -- 
    req_7798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(66), ack => array_obj_ref_3216_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Sample/ack
      -- 
    ack_7799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3216_index_offset_ack_0, ack => zeropad3D_E_CP_7148_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/array_obj_ref_3216_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_request/req
      -- 
    ack_7804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3216_index_offset_ack_1, ack => zeropad3D_E_CP_7148_elements(68)); -- 
    req_7813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(68), ack => addr_of_3217_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_request/ack
      -- 
    ack_7814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3217_final_reg_ack_0, ack => zeropad3D_E_CP_7148_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/addr_of_3217_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_word_addrgen/root_register_ack
      -- 
    ack_7819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3217_final_reg_ack_1, ack => zeropad3D_E_CP_7148_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/ptr_deref_3220_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/ptr_deref_3220_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/ptr_deref_3220_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/ptr_deref_3220_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/word_access_start/word_0/rr
      -- 
    rr_7857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(71), ack => ptr_deref_3220_store_0_req_0); -- 
    zeropad3D_E_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(64) & zeropad3D_E_CP_7148_elements(70);
      gj_zeropad3D_E_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Sample/word_access_start/word_0/ra
      -- 
    ra_7858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3220_store_0_ack_0, ack => zeropad3D_E_CP_7148_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/ptr_deref_3220_Update/word_access_complete/word_0/ca
      -- 
    ca_7869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3220_store_0_ack_1, ack => zeropad3D_E_CP_7148_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	111 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222__exit__
      -- CP-element group 74: 	 branch_block_stmt_2818/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_2818/assign_stmt_3122_to_assign_stmt_3222/$exit
      -- CP-element group 74: 	 branch_block_stmt_2818/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2818/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_E_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(59) & zeropad3D_E_CP_7148_elements(67) & zeropad3D_E_CP_7148_elements(73);
      gj_zeropad3D_E_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	111 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Sample/ra
      -- 
    ra_7881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3228_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	111 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243__entry__
      -- CP-element group 76: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242__exit__
      -- CP-element group 76: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/$exit
      -- CP-element group 76: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_2818/R_cmp145_3244_place
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_2818/if_stmt_3243_else_link/$entry
      -- 
    ca_7886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3228_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(76)); -- 
    branch_req_7894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(76), ack => if_stmt_3243_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	127 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187
      -- CP-element group 77: 	 branch_block_stmt_2818/assign_stmt_3255__exit__
      -- CP-element group 77: 	 branch_block_stmt_2818/assign_stmt_3255__entry__
      -- CP-element group 77: 	 branch_block_stmt_2818/merge_stmt_3249__exit__
      -- CP-element group 77: 	 branch_block_stmt_2818/if_stmt_3243_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_2818/if_stmt_3243_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xend_ifx_xthen147
      -- CP-element group 77: 	 branch_block_stmt_2818/assign_stmt_3255/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/assign_stmt_3255/$exit
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xend_ifx_xthen147_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xend_ifx_xthen147_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_2818/merge_stmt_3249_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_2818/merge_stmt_3249_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/merge_stmt_3249_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_2818/merge_stmt_3249_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3243_branch_ack_1, ack => zeropad3D_E_CP_7148_elements(77)); -- 
    rr_8256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(77), ack => type_cast_3323_inst_req_0); -- 
    cr_8261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(77), ack => type_cast_3323_inst_req_1); -- 
    rr_8279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(77), ack => type_cast_3317_inst_req_0); -- 
    cr_8284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(77), ack => type_cast_3317_inst_req_1); -- 
    rr_8302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(77), ack => type_cast_3310_inst_req_0); -- 
    cr_8307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(77), ack => type_cast_3310_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (24) 
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299__entry__
      -- CP-element group 78: 	 branch_block_stmt_2818/merge_stmt_3257__exit__
      -- CP-element group 78: 	 branch_block_stmt_2818/if_stmt_3243_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_2818/if_stmt_3243_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_2818/ifx_xend_ifx_xelse152
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_2818/ifx_xend_ifx_xelse152_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/ifx_xend_ifx_xelse152_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2818/merge_stmt_3257_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2818/merge_stmt_3257_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2818/merge_stmt_3257_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2818/merge_stmt_3257_PhiAck/dummy
      -- 
    else_choice_transition_7903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3243_branch_ack_0, ack => zeropad3D_E_CP_7148_elements(78)); -- 
    rr_7919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(78), ack => type_cast_3267_inst_req_0); -- 
    cr_7924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(78), ack => type_cast_3267_inst_req_1); -- 
    cr_7938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(78), ack => type_cast_3276_inst_req_1); -- 
    cr_7952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(78), ack => type_cast_3293_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Sample/ra
      -- 
    ra_7920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3267_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3267_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Sample/rr
      -- 
    ca_7925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3267_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(80)); -- 
    rr_7933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(80), ack => type_cast_3276_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Sample/ra
      -- 
    ra_7934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3276_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3276_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Sample/rr
      -- 
    ca_7939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3276_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(82)); -- 
    rr_7947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(82), ack => type_cast_3293_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Sample/ra
      -- 
    ra_7948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3293_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(83)); -- 
    -- CP-element group 84:  branch  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (13) 
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300__entry__
      -- CP-element group 84: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299__exit__
      -- CP-element group 84: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/$exit
      -- CP-element group 84: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_2818/assign_stmt_3263_to_assign_stmt_3299/type_cast_3293_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_2818/R_cmp179_3301_place
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_2818/if_stmt_3300_else_link/$entry
      -- 
    ca_7953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3293_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(84)); -- 
    branch_req_7961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(84), ack => if_stmt_3300_branch_req_0); -- 
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_2818/assign_stmt_3333__entry__
      -- CP-element group 85: 	 branch_block_stmt_2818/merge_stmt_3328__exit__
      -- CP-element group 85: 	 branch_block_stmt_2818/if_stmt_3300_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_2818/if_stmt_3300_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_2818/ifx_xelse152_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_2818/assign_stmt_3333/$entry
      -- CP-element group 85: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_2818/ifx_xelse152_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_2818/ifx_xelse152_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_2818/merge_stmt_3328_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_2818/merge_stmt_3328_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_2818/merge_stmt_3328_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_2818/merge_stmt_3328_PhiAck/dummy
      -- 
    if_choice_transition_7966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3300_branch_ack_1, ack => zeropad3D_E_CP_7148_elements(85)); -- 
    req_7983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(85), ack => WPIPE_Block4_complete_3330_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	115 
    -- CP-element group 86: 	116 
    -- CP-element group 86: 	118 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_2818/if_stmt_3300_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_2818/if_stmt_3300_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3307/$entry
      -- CP-element group 86: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/$entry
      -- 
    else_choice_transition_7970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3300_branch_ack_0, ack => zeropad3D_E_CP_7148_elements(86)); -- 
    rr_8199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(86), ack => type_cast_3325_inst_req_0); -- 
    cr_8204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(86), ack => type_cast_3325_inst_req_1); -- 
    rr_8222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(86), ack => type_cast_3319_inst_req_0); -- 
    cr_8227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(86), ack => type_cast_3319_inst_req_1); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_update_start_
      -- CP-element group 87: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Update/req
      -- 
    ack_7984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_complete_3330_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(87)); -- 
    req_7988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(87), ack => WPIPE_Block4_complete_3330_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_2818/$exit
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_2818/branch_block_stmt_2818__exit__
      -- CP-element group 88: 	 branch_block_stmt_2818/merge_stmt_3335__exit__
      -- CP-element group 88: 	 branch_block_stmt_2818/return__
      -- CP-element group 88: 	 branch_block_stmt_2818/assign_stmt_3333__exit__
      -- CP-element group 88: 	 branch_block_stmt_2818/assign_stmt_3333/$exit
      -- CP-element group 88: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_2818/assign_stmt_3333/WPIPE_Block4_complete_3330_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_2818/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_2818/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_2818/merge_stmt_3335_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_2818/merge_stmt_3335_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_2818/merge_stmt_3335_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_2818/merge_stmt_3335_PhiAck/dummy
      -- 
    ack_7989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block4_complete_3330_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(88)); -- 
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	94 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2965/$exit
      -- CP-element group 89: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2969_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_req
      -- 
    phi_stmt_2965_req_8000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2965_req_8000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(89), ack => phi_stmt_2965_req_0); -- 
    -- Element group zeropad3D_E_CP_7148_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_E_CP_7148_elements(32), ack => zeropad3D_E_CP_7148_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	32 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Sample/ra
      -- 
    ra_8017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2975_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/Update/ca
      -- 
    ca_8022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2975_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/$exit
      -- CP-element group 92: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/$exit
      -- CP-element group 92: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2975/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_req
      -- 
    phi_stmt_2972_req_8023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2972_req_8023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(92), ack => phi_stmt_2972_req_0); -- 
    zeropad3D_E_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(90) & zeropad3D_E_CP_7148_elements(91);
      gj_zeropad3D_E_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	32 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2978/$exit
      -- CP-element group 93: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2982_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_req
      -- 
    phi_stmt_2978_req_8031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2978_req_8031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(93), ack => phi_stmt_2978_req_0); -- 
    -- Element group zeropad3D_E_CP_7148_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => zeropad3D_E_CP_7148_elements(32), ack => zeropad3D_E_CP_7148_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	105 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2818/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_E_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(89) & zeropad3D_E_CP_7148_elements(92) & zeropad3D_E_CP_7148_elements(93);
      gj_zeropad3D_E_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Sample/ra
      -- 
    ra_8051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2971_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/Update/ca
      -- 
    ca_8056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2971_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/$exit
      -- CP-element group 97: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/$exit
      -- CP-element group 97: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_sources/type_cast_2971/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2965/phi_stmt_2965_req
      -- 
    phi_stmt_2965_req_8057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2965_req_8057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(97), ack => phi_stmt_2965_req_1); -- 
    zeropad3D_E_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_E_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(95) & zeropad3D_E_CP_7148_elements(96);
      gj_zeropad3D_E_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Sample/ra
      -- 
    ra_8074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2977_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/Update/ca
      -- 
    ca_8079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2977_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/$exit
      -- CP-element group 100: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/$exit
      -- CP-element group 100: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_sources/type_cast_2977/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2972/phi_stmt_2972_req
      -- 
    phi_stmt_2972_req_8080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2972_req_8080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(100), ack => phi_stmt_2972_req_1); -- 
    zeropad3D_E_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(98) & zeropad3D_E_CP_7148_elements(99);
      gj_zeropad3D_E_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Sample/ra
      -- 
    ra_8097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2984_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/Update/ca
      -- 
    ca_8102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2984_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/$exit
      -- CP-element group 103: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/$exit
      -- CP-element group 103: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_sources/type_cast_2984/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_2978/phi_stmt_2978_req
      -- 
    phi_stmt_2978_req_8103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2978_req_8103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(103), ack => phi_stmt_2978_req_1); -- 
    zeropad3D_E_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(101) & zeropad3D_E_CP_7148_elements(102);
      gj_zeropad3D_E_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_2818/ifx_xend187_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_E_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(97) & zeropad3D_E_CP_7148_elements(100) & zeropad3D_E_CP_7148_elements(103);
      gj_zeropad3D_E_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  merge  fork  transition  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	94 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2818/merge_stmt_2964_PhiReqMerge
      -- CP-element group 105: 	 branch_block_stmt_2818/merge_stmt_2964_PhiAck/$entry
      -- 
    zeropad3D_E_CP_7148_elements(105) <= OrReduce(zeropad3D_E_CP_7148_elements(94) & zeropad3D_E_CP_7148_elements(104));
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_2818/merge_stmt_2964_PhiAck/phi_stmt_2965_ack
      -- 
    phi_stmt_2965_ack_8108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2965_ack_0, ack => zeropad3D_E_CP_7148_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2818/merge_stmt_2964_PhiAck/phi_stmt_2972_ack
      -- 
    phi_stmt_2972_ack_8109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2972_ack_0, ack => zeropad3D_E_CP_7148_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2818/merge_stmt_2964_PhiAck/phi_stmt_2978_ack
      -- 
    phi_stmt_2978_ack_8110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2978_ack_0, ack => zeropad3D_E_CP_7148_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	33 
    -- CP-element group 109: 	34 
    -- CP-element group 109:  members (10) 
      -- CP-element group 109: 	 branch_block_stmt_2818/merge_stmt_2964__exit__
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015__entry__
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_update_start_
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/$entry
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_2818/assign_stmt_2990_to_assign_stmt_3015/type_cast_2989_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_2818/merge_stmt_2964_PhiAck/$exit
      -- 
    cr_7435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(109), ack => type_cast_2989_inst_req_1); -- 
    rr_7430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(109), ack => type_cast_2989_inst_req_0); -- 
    zeropad3D_E_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(106) & zeropad3D_E_CP_7148_elements(107) & zeropad3D_E_CP_7148_elements(108);
      gj_zeropad3D_E_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  merge  fork  transition  place  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	36 
    -- CP-element group 110: 	40 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	41 
    -- CP-element group 110: 	42 
    -- CP-element group 110: 	44 
    -- CP-element group 110: 	53 
    -- CP-element group 110: 	43 
    -- CP-element group 110: 	47 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	51 
    -- CP-element group 110:  members (33) 
      -- CP-element group 110: 	 branch_block_stmt_2818/merge_stmt_3059__exit__
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_update_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3063_update_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115__entry__
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3068_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_update_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/type_cast_3102_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_update_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_update_start
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/array_obj_ref_3108_final_index_sum_regn_Update/req
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/addr_of_3109_complete/req
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_update_start_
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/word_access_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/word_access_complete/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/assign_stmt_3064_to_assign_stmt_3115/ptr_deref_3112_Update/word_access_complete/word_0/cr
      -- CP-element group 110: 	 branch_block_stmt_2818/merge_stmt_3059_PhiReqMerge
      -- CP-element group 110: 	 branch_block_stmt_2818/merge_stmt_3059_PhiAck/$entry
      -- CP-element group 110: 	 branch_block_stmt_2818/merge_stmt_3059_PhiAck/$exit
      -- CP-element group 110: 	 branch_block_stmt_2818/merge_stmt_3059_PhiAck/dummy
      -- 
    rr_7502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => type_cast_3063_inst_req_0); -- 
    cr_7507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => type_cast_3063_inst_req_1); -- 
    rr_7516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => type_cast_3068_inst_req_0); -- 
    cr_7521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => type_cast_3068_inst_req_1); -- 
    cr_7535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => type_cast_3102_inst_req_1); -- 
    req_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => array_obj_ref_3108_index_offset_req_1); -- 
    req_7581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => addr_of_3109_final_reg_req_1); -- 
    cr_7631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(110), ack => ptr_deref_3112_store_0_req_1); -- 
    zeropad3D_E_CP_7148_elements(110) <= OrReduce(zeropad3D_E_CP_7148_elements(36) & zeropad3D_E_CP_7148_elements(40));
    -- CP-element group 111:  merge  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	54 
    -- CP-element group 111: 	74 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	75 
    -- CP-element group 111: 	76 
    -- CP-element group 111:  members (13) 
      -- CP-element group 111: 	 branch_block_stmt_2818/merge_stmt_3224__exit__
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242__entry__
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/$entry
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_update_start_
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_2818/assign_stmt_3229_to_assign_stmt_3242/type_cast_3228_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_2818/merge_stmt_3224_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_2818/merge_stmt_3224_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_2818/merge_stmt_3224_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_2818/merge_stmt_3224_PhiAck/dummy
      -- 
    rr_7880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(111), ack => type_cast_3228_inst_req_0); -- 
    cr_7885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(111), ack => type_cast_3228_inst_req_1); -- 
    zeropad3D_E_CP_7148_elements(111) <= OrReduce(zeropad3D_E_CP_7148_elements(54) & zeropad3D_E_CP_7148_elements(74));
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Sample/ra
      -- 
    ra_8200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3325_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/Update/ca
      -- 
    ca_8205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3325_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	119 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/$exit
      -- CP-element group 114: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/$exit
      -- CP-element group 114: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3325/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_req
      -- 
    phi_stmt_3320_req_8206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3320_req_8206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(114), ack => phi_stmt_3320_req_1); -- 
    zeropad3D_E_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(112) & zeropad3D_E_CP_7148_elements(113);
      gj_zeropad3D_E_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	86 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Sample/ra
      -- 
    ra_8223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3319_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/Update/ca
      -- 
    ca_8228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3319_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/$exit
      -- CP-element group 117: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/$exit
      -- CP-element group 117: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3319/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_req
      -- 
    phi_stmt_3314_req_8229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3314_req_8229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(117), ack => phi_stmt_3314_req_1); -- 
    zeropad3D_E_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(115) & zeropad3D_E_CP_7148_elements(116);
      gj_zeropad3D_E_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  output  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	86 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3307/$exit
      -- CP-element group 118: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3313_konst_delay_trans
      -- CP-element group 118: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_req
      -- 
    phi_stmt_3307_req_8237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3307_req_8237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(118), ack => phi_stmt_3307_req_1); -- 
    -- Element group zeropad3D_E_CP_7148_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => zeropad3D_E_CP_7148_elements(86), ack => zeropad3D_E_CP_7148_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  join  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	114 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	130 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_2818/ifx_xelse152_ifx_xend187_PhiReq/$exit
      -- 
    zeropad3D_E_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(114) & zeropad3D_E_CP_7148_elements(117) & zeropad3D_E_CP_7148_elements(118);
      gj_zeropad3D_E_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Sample/ra
      -- 
    ra_8257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3323_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/Update/ca
      -- 
    ca_8262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3323_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	129 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/$exit
      -- CP-element group 122: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/$exit
      -- CP-element group 122: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_sources/type_cast_3323/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3320/phi_stmt_3320_req
      -- 
    phi_stmt_3320_req_8263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3320_req_8263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(122), ack => phi_stmt_3320_req_0); -- 
    zeropad3D_E_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(120) & zeropad3D_E_CP_7148_elements(121);
      gj_zeropad3D_E_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Sample/ra
      -- 
    ra_8280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3317_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/Update/ca
      -- 
    ca_8285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3317_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/$exit
      -- CP-element group 125: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/$exit
      -- CP-element group 125: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_sources/type_cast_3317/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3314/phi_stmt_3314_req
      -- 
    phi_stmt_3314_req_8286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3314_req_8286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(125), ack => phi_stmt_3314_req_0); -- 
    zeropad3D_E_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(123) & zeropad3D_E_CP_7148_elements(124);
      gj_zeropad3D_E_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Sample/ra
      -- 
    ra_8303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3310_inst_ack_0, ack => zeropad3D_E_CP_7148_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	77 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/Update/ca
      -- 
    ca_8308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3310_inst_ack_1, ack => zeropad3D_E_CP_7148_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/$exit
      -- CP-element group 128: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/$exit
      -- CP-element group 128: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_sources/type_cast_3310/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/phi_stmt_3307/phi_stmt_3307_req
      -- 
    phi_stmt_3307_req_8309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3307_req_8309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_E_CP_7148_elements(128), ack => phi_stmt_3307_req_0); -- 
    zeropad3D_E_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(126) & zeropad3D_E_CP_7148_elements(127);
      gj_zeropad3D_E_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_2818/ifx_xthen147_ifx_xend187_PhiReq/$exit
      -- 
    zeropad3D_E_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(122) & zeropad3D_E_CP_7148_elements(125) & zeropad3D_E_CP_7148_elements(128);
      gj_zeropad3D_E_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_2818/merge_stmt_3306_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_2818/merge_stmt_3306_PhiAck/$entry
      -- 
    zeropad3D_E_CP_7148_elements(130) <= OrReduce(zeropad3D_E_CP_7148_elements(119) & zeropad3D_E_CP_7148_elements(129));
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_2818/merge_stmt_3306_PhiAck/phi_stmt_3307_ack
      -- 
    phi_stmt_3307_ack_8314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3307_ack_0, ack => zeropad3D_E_CP_7148_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_2818/merge_stmt_3306_PhiAck/phi_stmt_3314_ack
      -- 
    phi_stmt_3314_ack_8315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3314_ack_0, ack => zeropad3D_E_CP_7148_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_2818/merge_stmt_3306_PhiAck/phi_stmt_3320_ack
      -- 
    phi_stmt_3320_ack_8316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3320_ack_0, ack => zeropad3D_E_CP_7148_elements(133)); -- 
    -- CP-element group 134:  join  transition  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	1 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_2818/merge_stmt_3306_PhiAck/$exit
      -- 
    zeropad3D_E_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_E_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_E_CP_7148_elements(131) & zeropad3D_E_CP_7148_elements(132) & zeropad3D_E_CP_7148_elements(133);
      gj_zeropad3D_E_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_E_CP_7148_elements(134), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2892_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2960_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3096_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3179_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3204_wire : std_logic_vector(31 downto 0);
    signal R_idxprom132_3190_resized : std_logic_vector(13 downto 0);
    signal R_idxprom132_3190_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom137_3215_resized : std_logic_vector(13 downto 0);
    signal R_idxprom137_3215_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3107_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3107_scaled : std_logic_vector(13 downto 0);
    signal add104_3147 : std_logic_vector(31 downto 0);
    signal add113_3152 : std_logic_vector(31 downto 0);
    signal add123_3167 : std_logic_vector(31 downto 0);
    signal add129_3172 : std_logic_vector(31 downto 0);
    signal add142_3235 : std_logic_vector(31 downto 0);
    signal add150_3255 : std_logic_vector(15 downto 0);
    signal add161_2911 : std_logic_vector(31 downto 0);
    signal add178_2932 : std_logic_vector(31 downto 0);
    signal add75_2942 : std_logic_vector(31 downto 0);
    signal add86_3084 : std_logic_vector(31 downto 0);
    signal add92_3089 : std_logic_vector(31 downto 0);
    signal add_2937 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3108_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3108_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3108_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3108_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3108_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3108_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3191_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3191_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3191_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3191_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3191_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3191_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3216_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3216_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3216_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3216_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3216_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3216_root_address : std_logic_vector(13 downto 0);
    signal arrayidx133_3193 : std_logic_vector(31 downto 0);
    signal arrayidx138_3218 : std_logic_vector(31 downto 0);
    signal arrayidx_3110 : std_logic_vector(31 downto 0);
    signal call1_2824 : std_logic_vector(7 downto 0);
    signal call2_2827 : std_logic_vector(7 downto 0);
    signal call3_2830 : std_logic_vector(7 downto 0);
    signal call4_2833 : std_logic_vector(7 downto 0);
    signal call5_2836 : std_logic_vector(7 downto 0);
    signal call6_2839 : std_logic_vector(7 downto 0);
    signal call_2821 : std_logic_vector(7 downto 0);
    signal cmp145_3242 : std_logic_vector(0 downto 0);
    signal cmp162_3273 : std_logic_vector(0 downto 0);
    signal cmp179_3299 : std_logic_vector(0 downto 0);
    signal cmp58_3010 : std_logic_vector(0 downto 0);
    signal cmp65_3034 : std_logic_vector(0 downto 0);
    signal cmp65x_xnot_3040 : std_logic_vector(0 downto 0);
    signal cmp76_3047 : std_logic_vector(0 downto 0);
    signal cmp_2997 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_3003 : std_logic_vector(0 downto 0);
    signal conv106_2962 : std_logic_vector(31 downto 0);
    signal conv141_3229 : std_logic_vector(31 downto 0);
    signal conv155_3268 : std_logic_vector(31 downto 0);
    signal conv170_3294 : std_logic_vector(31 downto 0);
    signal conv172_2915 : std_logic_vector(31 downto 0);
    signal conv31_2854 : std_logic_vector(31 downto 0);
    signal conv33_2858 : std_logic_vector(31 downto 0);
    signal conv37_2862 : std_logic_vector(31 downto 0);
    signal conv39_2866 : std_logic_vector(31 downto 0);
    signal conv46_2990 : std_logic_vector(31 downto 0);
    signal conv48_2875 : std_logic_vector(31 downto 0);
    signal conv62_3027 : std_logic_vector(31 downto 0);
    signal conv80_3064 : std_logic_vector(31 downto 0);
    signal conv82_2879 : std_logic_vector(31 downto 0);
    signal conv84_3069 : std_logic_vector(31 downto 0);
    signal conv88_2894 : std_logic_vector(31 downto 0);
    signal conv96_3122 : std_logic_vector(31 downto 0);
    signal conv_2844 : std_logic_vector(15 downto 0);
    signal div158_2900 : std_logic_vector(31 downto 0);
    signal div174_2927 : std_logic_vector(31 downto 0);
    signal div_2850 : std_logic_vector(15 downto 0);
    signal idxprom132_3186 : std_logic_vector(63 downto 0);
    signal idxprom137_3211 : std_logic_vector(63 downto 0);
    signal idxprom_3103 : std_logic_vector(63 downto 0);
    signal inc167_3277 : std_logic_vector(15 downto 0);
    signal inc167x_xix_x2_3282 : std_logic_vector(15 downto 0);
    signal inc_3263 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_3314 : std_logic_vector(15 downto 0);
    signal ix_x2_2972 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_3320 : std_logic_vector(15 downto 0);
    signal jx_x1_2978 : std_logic_vector(15 downto 0);
    signal jx_x2_3289 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_3307 : std_logic_vector(15 downto 0);
    signal kx_x1_2965 : std_logic_vector(15 downto 0);
    signal mul103_3132 : std_logic_vector(31 downto 0);
    signal mul112_3142 : std_logic_vector(31 downto 0);
    signal mul122_3157 : std_logic_vector(31 downto 0);
    signal mul128_3162 : std_logic_vector(31 downto 0);
    signal mul173_2921 : std_logic_vector(31 downto 0);
    signal mul40_2871 : std_logic_vector(31 downto 0);
    signal mul85_3074 : std_logic_vector(31 downto 0);
    signal mul91_3079 : std_logic_vector(31 downto 0);
    signal mul_2948 : std_logic_vector(31 downto 0);
    signal orx_xcond193_3052 : std_logic_vector(0 downto 0);
    signal orx_xcond_3015 : std_logic_vector(0 downto 0);
    signal ptr_deref_3112_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3112_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3112_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3112_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3112_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3112_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3196_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3196_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3220_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3220_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3220_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3220_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3220_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3220_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext192_2885 : std_logic_vector(31 downto 0);
    signal sext_2953 : std_logic_vector(31 downto 0);
    signal shl_2906 : std_logic_vector(31 downto 0);
    signal shr131_3181 : std_logic_vector(31 downto 0);
    signal shr136_3206 : std_logic_vector(31 downto 0);
    signal shr_3098 : std_logic_vector(31 downto 0);
    signal sub111_3137 : std_logic_vector(31 downto 0);
    signal sub_3127 : std_logic_vector(31 downto 0);
    signal tmp134_3197 : std_logic_vector(63 downto 0);
    signal type_cast_2848_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2883_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2888_wire : std_logic_vector(31 downto 0);
    signal type_cast_2891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2904_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2919_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2925_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2946_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2956_wire : std_logic_vector(31 downto 0);
    signal type_cast_2959_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2969_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2971_wire : std_logic_vector(15 downto 0);
    signal type_cast_2975_wire : std_logic_vector(15 downto 0);
    signal type_cast_2977_wire : std_logic_vector(15 downto 0);
    signal type_cast_2982_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2984_wire : std_logic_vector(15 downto 0);
    signal type_cast_2988_wire : std_logic_vector(31 downto 0);
    signal type_cast_2993_wire : std_logic_vector(31 downto 0);
    signal type_cast_2995_wire : std_logic_vector(31 downto 0);
    signal type_cast_3001_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3006_wire : std_logic_vector(31 downto 0);
    signal type_cast_3008_wire : std_logic_vector(31 downto 0);
    signal type_cast_3025_wire : std_logic_vector(31 downto 0);
    signal type_cast_3030_wire : std_logic_vector(31 downto 0);
    signal type_cast_3032_wire : std_logic_vector(31 downto 0);
    signal type_cast_3038_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3043_wire : std_logic_vector(31 downto 0);
    signal type_cast_3045_wire : std_logic_vector(31 downto 0);
    signal type_cast_3062_wire : std_logic_vector(31 downto 0);
    signal type_cast_3067_wire : std_logic_vector(31 downto 0);
    signal type_cast_3092_wire : std_logic_vector(31 downto 0);
    signal type_cast_3095_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3101_wire : std_logic_vector(63 downto 0);
    signal type_cast_3114_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3120_wire : std_logic_vector(31 downto 0);
    signal type_cast_3175_wire : std_logic_vector(31 downto 0);
    signal type_cast_3178_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3184_wire : std_logic_vector(63 downto 0);
    signal type_cast_3200_wire : std_logic_vector(31 downto 0);
    signal type_cast_3203_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3209_wire : std_logic_vector(63 downto 0);
    signal type_cast_3227_wire : std_logic_vector(31 downto 0);
    signal type_cast_3233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3238_wire : std_logic_vector(31 downto 0);
    signal type_cast_3240_wire : std_logic_vector(31 downto 0);
    signal type_cast_3253_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3261_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3266_wire : std_logic_vector(31 downto 0);
    signal type_cast_3286_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3292_wire : std_logic_vector(31 downto 0);
    signal type_cast_3310_wire : std_logic_vector(15 downto 0);
    signal type_cast_3313_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3317_wire : std_logic_vector(15 downto 0);
    signal type_cast_3319_wire : std_logic_vector(15 downto 0);
    signal type_cast_3323_wire : std_logic_vector(15 downto 0);
    signal type_cast_3325_wire : std_logic_vector(15 downto 0);
    signal type_cast_3332_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_3108_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3108_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3108_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3108_resized_base_address <= "00000000000000";
    array_obj_ref_3191_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3191_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3191_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3191_resized_base_address <= "00000000000000";
    array_obj_ref_3216_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3216_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3216_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3216_resized_base_address <= "00000000000000";
    ptr_deref_3112_word_offset_0 <= "00000000000000";
    ptr_deref_3196_word_offset_0 <= "00000000000000";
    ptr_deref_3220_word_offset_0 <= "00000000000000";
    type_cast_2848_wire_constant <= "0000000000000001";
    type_cast_2883_wire_constant <= "00000000000000000000000000010000";
    type_cast_2891_wire_constant <= "00000000000000000000000000010000";
    type_cast_2898_wire_constant <= "00000000000000000000000000000001";
    type_cast_2904_wire_constant <= "00000000000000000000000000000001";
    type_cast_2919_wire_constant <= "00000000000000000000000000000011";
    type_cast_2925_wire_constant <= "00000000000000000000000000000010";
    type_cast_2946_wire_constant <= "00000000000000000000000000010000";
    type_cast_2959_wire_constant <= "00000000000000000000000000010000";
    type_cast_2969_wire_constant <= "0000000000000000";
    type_cast_2982_wire_constant <= "0000000000000000";
    type_cast_3001_wire_constant <= "1";
    type_cast_3038_wire_constant <= "1";
    type_cast_3095_wire_constant <= "00000000000000000000000000000010";
    type_cast_3114_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3178_wire_constant <= "00000000000000000000000000000010";
    type_cast_3203_wire_constant <= "00000000000000000000000000000010";
    type_cast_3233_wire_constant <= "00000000000000000000000000000100";
    type_cast_3253_wire_constant <= "0000000000000100";
    type_cast_3261_wire_constant <= "0000000000000001";
    type_cast_3286_wire_constant <= "0000000000000000";
    type_cast_3313_wire_constant <= "0000000000000000";
    type_cast_3332_wire_constant <= "00000001";
    phi_stmt_2965: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2969_wire_constant & type_cast_2971_wire;
      req <= phi_stmt_2965_req_0 & phi_stmt_2965_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2965",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2965_ack_0,
          idata => idata,
          odata => kx_x1_2965,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2965
    phi_stmt_2972: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2975_wire & type_cast_2977_wire;
      req <= phi_stmt_2972_req_0 & phi_stmt_2972_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2972",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2972_ack_0,
          idata => idata,
          odata => ix_x2_2972,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2972
    phi_stmt_2978: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2982_wire_constant & type_cast_2984_wire;
      req <= phi_stmt_2978_req_0 & phi_stmt_2978_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2978",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2978_ack_0,
          idata => idata,
          odata => jx_x1_2978,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2978
    phi_stmt_3307: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3310_wire & type_cast_3313_wire_constant;
      req <= phi_stmt_3307_req_0 & phi_stmt_3307_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3307",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3307_ack_0,
          idata => idata,
          odata => kx_x0x_xph_3307,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3307
    phi_stmt_3314: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3317_wire & type_cast_3319_wire;
      req <= phi_stmt_3314_req_0 & phi_stmt_3314_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3314",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3314_ack_0,
          idata => idata,
          odata => ix_x1x_xph_3314,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3314
    phi_stmt_3320: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3323_wire & type_cast_3325_wire;
      req <= phi_stmt_3320_req_0 & phi_stmt_3320_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3320",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3320_ack_0,
          idata => idata,
          odata => jx_x0x_xph_3320,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3320
    -- flow-through select operator MUX_3288_inst
    jx_x2_3289 <= type_cast_3286_wire_constant when (cmp162_3273(0) /=  '0') else inc_3263;
    addr_of_3109_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3109_final_reg_req_0;
      addr_of_3109_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3109_final_reg_req_1;
      addr_of_3109_final_reg_ack_1<= rack(0);
      addr_of_3109_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3109_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3108_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3192_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3192_final_reg_req_0;
      addr_of_3192_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3192_final_reg_req_1;
      addr_of_3192_final_reg_ack_1<= rack(0);
      addr_of_3192_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3192_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3191_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx133_3193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3217_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3217_final_reg_req_0;
      addr_of_3217_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3217_final_reg_req_1;
      addr_of_3217_final_reg_ack_1<= rack(0);
      addr_of_3217_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3217_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3216_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx138_3218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2843_inst_req_0;
      type_cast_2843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2843_inst_req_1;
      type_cast_2843_inst_ack_1<= rack(0);
      type_cast_2843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2853_inst_req_0;
      type_cast_2853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2853_inst_req_1;
      type_cast_2853_inst_ack_1<= rack(0);
      type_cast_2853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_2827,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_2854,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2857_inst_req_0;
      type_cast_2857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2857_inst_req_1;
      type_cast_2857_inst_ack_1<= rack(0);
      type_cast_2857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_2858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2861_inst_req_0;
      type_cast_2861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2861_inst_req_1;
      type_cast_2861_inst_ack_1<= rack(0);
      type_cast_2861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_2836,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_2862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2865_inst_req_0;
      type_cast_2865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2865_inst_req_1;
      type_cast_2865_inst_ack_1<= rack(0);
      type_cast_2865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_2833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_2866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2874_inst_req_0;
      type_cast_2874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2874_inst_req_1;
      type_cast_2874_inst_ack_1<= rack(0);
      type_cast_2874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_2839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_2875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2878_inst_req_0;
      type_cast_2878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2878_inst_req_1;
      type_cast_2878_inst_ack_1<= rack(0);
      type_cast_2878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2878_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_2836,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_2879,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2888_inst
    process(sext192_2885) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext192_2885(31 downto 0);
      type_cast_2888_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2893_inst
    process(ASHR_i32_i32_2892_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2892_wire(31 downto 0);
      conv88_2894 <= tmp_var; -- 
    end process;
    type_cast_2914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2914_inst_req_0;
      type_cast_2914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2914_inst_req_1;
      type_cast_2914_inst_ack_1<= rack(0);
      type_cast_2914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv172_2915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2956_inst
    process(sext_2953) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2953(31 downto 0);
      type_cast_2956_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2961_inst
    process(ASHR_i32_i32_2960_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2960_wire(31 downto 0);
      conv106_2962 <= tmp_var; -- 
    end process;
    type_cast_2971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2971_inst_req_0;
      type_cast_2971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2971_inst_req_1;
      type_cast_2971_inst_ack_1<= rack(0);
      type_cast_2971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_3307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2971_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2975_inst_req_0;
      type_cast_2975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2975_inst_req_1;
      type_cast_2975_inst_ack_1<= rack(0);
      type_cast_2975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2975_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2977_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2977_inst_req_0;
      type_cast_2977_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2977_inst_req_1;
      type_cast_2977_inst_ack_1<= rack(0);
      type_cast_2977_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2977_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_3314,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2977_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2984_inst_req_0;
      type_cast_2984_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2984_inst_req_1;
      type_cast_2984_inst_ack_1<= rack(0);
      type_cast_2984_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_3320,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2984_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2989_inst_req_0;
      type_cast_2989_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2989_inst_req_1;
      type_cast_2989_inst_ack_1<= rack(0);
      type_cast_2989_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2989_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2988_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_2990,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2993_inst
    process(conv46_2990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_2990(31 downto 0);
      type_cast_2993_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2995_inst
    process(conv48_2875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_2875(31 downto 0);
      type_cast_2995_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3006_inst
    process(conv46_2990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_2990(31 downto 0);
      type_cast_3006_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3008_inst
    process(add_2937) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_2937(31 downto 0);
      type_cast_3008_wire <= tmp_var; -- 
    end process;
    type_cast_3026_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3026_inst_req_0;
      type_cast_3026_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3026_inst_req_1;
      type_cast_3026_inst_ack_1<= rack(0);
      type_cast_3026_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3026_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3025_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_3027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3030_inst
    process(conv62_3027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv62_3027(31 downto 0);
      type_cast_3030_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3032_inst
    process(conv48_2875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_2875(31 downto 0);
      type_cast_3032_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3043_inst
    process(conv62_3027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv62_3027(31 downto 0);
      type_cast_3043_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3045_inst
    process(add75_2942) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add75_2942(31 downto 0);
      type_cast_3045_wire <= tmp_var; -- 
    end process;
    type_cast_3063_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3063_inst_req_0;
      type_cast_3063_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3063_inst_req_1;
      type_cast_3063_inst_ack_1<= rack(0);
      type_cast_3063_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3063_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3062_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_3064,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3068_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3068_inst_req_0;
      type_cast_3068_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3068_inst_req_1;
      type_cast_3068_inst_ack_1<= rack(0);
      type_cast_3068_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3068_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3067_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_3069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3092_inst
    process(add92_3089) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add92_3089(31 downto 0);
      type_cast_3092_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3097_inst
    process(ASHR_i32_i32_3096_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3096_wire(31 downto 0);
      shr_3098 <= tmp_var; -- 
    end process;
    type_cast_3102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3102_inst_req_0;
      type_cast_3102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3102_inst_req_1;
      type_cast_3102_inst_ack_1<= rack(0);
      type_cast_3102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3101_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3121_inst_req_0;
      type_cast_3121_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3121_inst_req_1;
      type_cast_3121_inst_ack_1<= rack(0);
      type_cast_3121_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3121_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3120_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_3122,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3175_inst
    process(add113_3152) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add113_3152(31 downto 0);
      type_cast_3175_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3180_inst
    process(ASHR_i32_i32_3179_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3179_wire(31 downto 0);
      shr131_3181 <= tmp_var; -- 
    end process;
    type_cast_3185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3185_inst_req_0;
      type_cast_3185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3185_inst_req_1;
      type_cast_3185_inst_ack_1<= rack(0);
      type_cast_3185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3184_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom132_3186,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3200_inst
    process(add129_3172) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add129_3172(31 downto 0);
      type_cast_3200_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3205_inst
    process(ASHR_i32_i32_3204_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3204_wire(31 downto 0);
      shr136_3206 <= tmp_var; -- 
    end process;
    type_cast_3210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3210_inst_req_0;
      type_cast_3210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3210_inst_req_1;
      type_cast_3210_inst_ack_1<= rack(0);
      type_cast_3210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3209_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom137_3211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3228_inst_req_0;
      type_cast_3228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3228_inst_req_1;
      type_cast_3228_inst_ack_1<= rack(0);
      type_cast_3228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3227_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_3229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3238_inst
    process(add142_3235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add142_3235(31 downto 0);
      type_cast_3238_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3240_inst
    process(conv31_2854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv31_2854(31 downto 0);
      type_cast_3240_wire <= tmp_var; -- 
    end process;
    type_cast_3267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3267_inst_req_0;
      type_cast_3267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3267_inst_req_1;
      type_cast_3267_inst_ack_1<= rack(0);
      type_cast_3267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3266_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_3268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3276_inst_req_0;
      type_cast_3276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3276_inst_req_1;
      type_cast_3276_inst_ack_1<= rack(0);
      type_cast_3276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp162_3273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc167_3277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3293_inst_req_0;
      type_cast_3293_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3293_inst_req_1;
      type_cast_3293_inst_ack_1<= rack(0);
      type_cast_3293_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3293_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3292_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_3294,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3310_inst_req_0;
      type_cast_3310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3310_inst_req_1;
      type_cast_3310_inst_ack_1<= rack(0);
      type_cast_3310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add150_3255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3310_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3317_inst_req_0;
      type_cast_3317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3317_inst_req_1;
      type_cast_3317_inst_ack_1<= rack(0);
      type_cast_3317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_2972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3317_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3319_inst_req_0;
      type_cast_3319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3319_inst_req_1;
      type_cast_3319_inst_ack_1<= rack(0);
      type_cast_3319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc167x_xix_x2_3282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3319_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3323_inst_req_0;
      type_cast_3323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3323_inst_req_1;
      type_cast_3323_inst_ack_1<= rack(0);
      type_cast_3323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_2978,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3323_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3325_inst_req_0;
      type_cast_3325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3325_inst_req_1;
      type_cast_3325_inst_ack_1<= rack(0);
      type_cast_3325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_3289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3325_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_3108_index_1_rename
    process(R_idxprom_3107_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3107_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3107_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3108_index_1_resize
    process(idxprom_3103) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3103;
      ov := iv(13 downto 0);
      R_idxprom_3107_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3108_root_address_inst
    process(array_obj_ref_3108_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3108_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3108_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3191_index_1_rename
    process(R_idxprom132_3190_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom132_3190_resized;
      ov(13 downto 0) := iv;
      R_idxprom132_3190_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3191_index_1_resize
    process(idxprom132_3186) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom132_3186;
      ov := iv(13 downto 0);
      R_idxprom132_3190_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3191_root_address_inst
    process(array_obj_ref_3191_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3191_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3191_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3216_index_1_rename
    process(R_idxprom137_3215_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom137_3215_resized;
      ov(13 downto 0) := iv;
      R_idxprom137_3215_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3216_index_1_resize
    process(idxprom137_3211) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom137_3211;
      ov := iv(13 downto 0);
      R_idxprom137_3215_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3216_root_address_inst
    process(array_obj_ref_3216_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3216_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3216_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3112_addr_0
    process(ptr_deref_3112_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3112_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3112_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3112_base_resize
    process(arrayidx_3110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3110;
      ov := iv(13 downto 0);
      ptr_deref_3112_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3112_gather_scatter
    process(type_cast_3114_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3114_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3112_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3112_root_address_inst
    process(ptr_deref_3112_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3112_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3112_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_addr_0
    process(ptr_deref_3196_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3196_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3196_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_base_resize
    process(arrayidx133_3193) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx133_3193;
      ov := iv(13 downto 0);
      ptr_deref_3196_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_gather_scatter
    process(ptr_deref_3196_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3196_data_0;
      ov(63 downto 0) := iv;
      tmp134_3197 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3196_root_address_inst
    process(ptr_deref_3196_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3196_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3196_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3220_addr_0
    process(ptr_deref_3220_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3220_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3220_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3220_base_resize
    process(arrayidx138_3218) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx138_3218;
      ov := iv(13 downto 0);
      ptr_deref_3220_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3220_gather_scatter
    process(tmp134_3197) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp134_3197;
      ov(63 downto 0) := iv;
      ptr_deref_3220_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3220_root_address_inst
    process(ptr_deref_3220_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3220_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3220_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3016_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_3015;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3016_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3016_branch_req_0,
          ack0 => if_stmt_3016_branch_ack_0,
          ack1 => if_stmt_3016_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3053_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond193_3052;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3053_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3053_branch_req_0,
          ack0 => if_stmt_3053_branch_ack_0,
          ack1 => if_stmt_3053_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3243_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp145_3242;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3243_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3243_branch_req_0,
          ack0 => if_stmt_3243_branch_ack_0,
          ack1 => if_stmt_3243_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3300_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp179_3299;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3300_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3300_branch_req_0,
          ack0 => if_stmt_3300_branch_ack_0,
          ack1 => if_stmt_3300_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3254_inst
    process(kx_x1_2965) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_2965, type_cast_3253_wire_constant, tmp_var);
      add150_3255 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3262_inst
    process(jx_x1_2978) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_2978, type_cast_3261_wire_constant, tmp_var);
      inc_3263 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3281_inst
    process(inc167_3277, ix_x2_2972) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc167_3277, ix_x2_2972, tmp_var);
      inc167x_xix_x2_3282 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2910_inst
    process(shl_2906, div158_2900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_2906, div158_2900, tmp_var);
      add161_2911 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2931_inst
    process(shl_2906, div174_2927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_2906, div174_2927, tmp_var);
      add178_2932 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2936_inst
    process(conv48_2875, div174_2927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv48_2875, div174_2927, tmp_var);
      add_2937 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2941_inst
    process(conv48_2875, div158_2900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv48_2875, div158_2900, tmp_var);
      add75_2942 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3083_inst
    process(mul91_3079, conv80_3064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul91_3079, conv80_3064, tmp_var);
      add86_3084 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3088_inst
    process(add86_3084, mul85_3074) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add86_3084, mul85_3074, tmp_var);
      add92_3089 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3146_inst
    process(mul112_3142, conv96_3122) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul112_3142, conv96_3122, tmp_var);
      add104_3147 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3151_inst
    process(add104_3147, mul103_3132) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add104_3147, mul103_3132, tmp_var);
      add113_3152 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3166_inst
    process(mul128_3162, conv96_3122) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul128_3162, conv96_3122, tmp_var);
      add123_3167 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3171_inst
    process(add123_3167, mul122_3157) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add123_3167, mul122_3157, tmp_var);
      add129_3172 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3234_inst
    process(conv141_3229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv141_3229, type_cast_3233_wire_constant, tmp_var);
      add142_3235 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3014_inst
    process(cmpx_xnot_3003, cmp58_3010) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_3003, cmp58_3010, tmp_var);
      orx_xcond_3015 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3051_inst
    process(cmp65x_xnot_3040, cmp76_3047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp65x_xnot_3040, cmp76_3047, tmp_var);
      orx_xcond193_3052 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2892_inst
    process(type_cast_2888_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2888_wire, type_cast_2891_wire_constant, tmp_var);
      ASHR_i32_i32_2892_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2960_inst
    process(type_cast_2956_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2956_wire, type_cast_2959_wire_constant, tmp_var);
      ASHR_i32_i32_2960_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3096_inst
    process(type_cast_3092_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3092_wire, type_cast_3095_wire_constant, tmp_var);
      ASHR_i32_i32_3096_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3179_inst
    process(type_cast_3175_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3175_wire, type_cast_3178_wire_constant, tmp_var);
      ASHR_i32_i32_3179_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3204_inst
    process(type_cast_3200_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3200_wire, type_cast_3203_wire_constant, tmp_var);
      ASHR_i32_i32_3204_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3272_inst
    process(conv155_3268, add161_2911) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv155_3268, add161_2911, tmp_var);
      cmp162_3273 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3298_inst
    process(conv170_3294, add178_2932) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv170_3294, add178_2932, tmp_var);
      cmp179_3299 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2849_inst
    process(conv_2844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_2844, type_cast_2848_wire_constant, tmp_var);
      div_2850 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2899_inst
    process(conv33_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv33_2858, type_cast_2898_wire_constant, tmp_var);
      div158_2900 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2926_inst
    process(mul173_2921) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul173_2921, type_cast_2925_wire_constant, tmp_var);
      div174_2927 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2870_inst
    process(conv37_2862, conv39_2866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_2862, conv39_2866, tmp_var);
      mul40_2871 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2920_inst
    process(conv172_2915) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv172_2915, type_cast_2919_wire_constant, tmp_var);
      mul173_2921 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2952_inst
    process(mul_2948, conv31_2854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_2948, conv31_2854, tmp_var);
      sext_2953 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3073_inst
    process(conv84_3069, conv82_2879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_3069, conv82_2879, tmp_var);
      mul85_3074 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3078_inst
    process(conv46_2990, conv88_2894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_2990, conv88_2894, tmp_var);
      mul91_3079 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3131_inst
    process(sub_3127, conv31_2854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_3127, conv31_2854, tmp_var);
      mul103_3132 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3141_inst
    process(sub111_3137, conv106_2962) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub111_3137, conv106_2962, tmp_var);
      mul112_3142 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3156_inst
    process(conv62_3027, conv82_2879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv62_3027, conv82_2879, tmp_var);
      mul122_3157 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3161_inst
    process(conv46_2990, conv88_2894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_2990, conv88_2894, tmp_var);
      mul128_3162 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2884_inst
    process(mul40_2871) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul40_2871, type_cast_2883_wire_constant, tmp_var);
      sext192_2885 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2905_inst
    process(conv48_2875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_2875, type_cast_2904_wire_constant, tmp_var);
      shl_2906 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2947_inst
    process(conv33_2858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv33_2858, type_cast_2946_wire_constant, tmp_var);
      mul_2948 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2996_inst
    process(type_cast_2993_wire, type_cast_2995_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2993_wire, type_cast_2995_wire, tmp_var);
      cmp_2997 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3009_inst
    process(type_cast_3006_wire, type_cast_3008_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3006_wire, type_cast_3008_wire, tmp_var);
      cmp58_3010 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3033_inst
    process(type_cast_3030_wire, type_cast_3032_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3030_wire, type_cast_3032_wire, tmp_var);
      cmp65_3034 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3046_inst
    process(type_cast_3043_wire, type_cast_3045_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3043_wire, type_cast_3045_wire, tmp_var);
      cmp76_3047 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3241_inst
    process(type_cast_3238_wire, type_cast_3240_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3238_wire, type_cast_3240_wire, tmp_var);
      cmp145_3242 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3126_inst
    process(conv62_3027, conv48_2875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv62_3027, conv48_2875, tmp_var);
      sub_3127 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3136_inst
    process(conv46_2990, conv48_2875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv46_2990, conv48_2875, tmp_var);
      sub111_3137 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3002_inst
    process(cmp_2997) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_2997, type_cast_3001_wire_constant, tmp_var);
      cmpx_xnot_3003 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3039_inst
    process(cmp65_3034) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp65_3034, type_cast_3038_wire_constant, tmp_var);
      cmp65x_xnot_3040 <= tmp_var; --
    end process;
    -- shared split operator group (47) : array_obj_ref_3108_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3107_scaled;
      array_obj_ref_3108_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3108_index_offset_req_0;
      array_obj_ref_3108_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3108_index_offset_req_1;
      array_obj_ref_3108_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_3191_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom132_3190_scaled;
      array_obj_ref_3191_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3191_index_offset_req_0;
      array_obj_ref_3191_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3191_index_offset_req_1;
      array_obj_ref_3191_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : array_obj_ref_3216_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom137_3215_scaled;
      array_obj_ref_3216_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3216_index_offset_req_0;
      array_obj_ref_3216_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3216_index_offset_req_1;
      array_obj_ref_3216_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- unary operator type_cast_2988_inst
    process(ix_x2_2972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_2972, tmp_var);
      type_cast_2988_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3025_inst
    process(jx_x1_2978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2978, tmp_var);
      type_cast_3025_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3062_inst
    process(kx_x1_2965) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2965, tmp_var);
      type_cast_3062_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3067_inst
    process(jx_x1_2978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2978, tmp_var);
      type_cast_3067_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3101_inst
    process(shr_3098) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3098, tmp_var);
      type_cast_3101_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3120_inst
    process(kx_x1_2965) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2965, tmp_var);
      type_cast_3120_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3184_inst
    process(shr131_3181) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr131_3181, tmp_var);
      type_cast_3184_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3209_inst
    process(shr136_3206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr136_3206, tmp_var);
      type_cast_3209_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3227_inst
    process(kx_x1_2965) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2965, tmp_var);
      type_cast_3227_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3266_inst
    process(inc_3263) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3263, tmp_var);
      type_cast_3266_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3292_inst
    process(inc167x_xix_x2_3282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc167x_xix_x2_3282, tmp_var);
      type_cast_3292_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_3196_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3196_load_0_req_0;
      ptr_deref_3196_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3196_load_0_req_1;
      ptr_deref_3196_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3196_word_address_0;
      ptr_deref_3196_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3112_store_0 ptr_deref_3220_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3112_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3220_store_0_req_0;
      ptr_deref_3112_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3220_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3112_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3220_store_0_req_1;
      ptr_deref_3112_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3220_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3112_word_address_0 & ptr_deref_3220_word_address_0;
      data_in <= ptr_deref_3112_data_0 & ptr_deref_3220_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block4_starting_2838_inst RPIPE_Block4_starting_2835_inst RPIPE_Block4_starting_2832_inst RPIPE_Block4_starting_2829_inst RPIPE_Block4_starting_2826_inst RPIPE_Block4_starting_2823_inst RPIPE_Block4_starting_2820_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block4_starting_2838_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block4_starting_2835_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block4_starting_2832_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block4_starting_2829_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block4_starting_2826_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block4_starting_2823_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block4_starting_2820_inst_req_0;
      RPIPE_Block4_starting_2838_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block4_starting_2835_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block4_starting_2832_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block4_starting_2829_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block4_starting_2826_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block4_starting_2823_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block4_starting_2820_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block4_starting_2838_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block4_starting_2835_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block4_starting_2832_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block4_starting_2829_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block4_starting_2826_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block4_starting_2823_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block4_starting_2820_inst_req_1;
      RPIPE_Block4_starting_2838_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block4_starting_2835_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block4_starting_2832_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block4_starting_2829_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block4_starting_2826_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block4_starting_2823_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block4_starting_2820_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call6_2839 <= data_out(55 downto 48);
      call5_2836 <= data_out(47 downto 40);
      call4_2833 <= data_out(39 downto 32);
      call3_2830 <= data_out(31 downto 24);
      call2_2827 <= data_out(23 downto 16);
      call1_2824 <= data_out(15 downto 8);
      call_2821 <= data_out(7 downto 0);
      Block4_starting_read_0_gI: SplitGuardInterface generic map(name => "Block4_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block4_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block4_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block4_starting_pipe_read_req(0),
          oack => Block4_starting_pipe_read_ack(0),
          odata => Block4_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block4_complete_3330_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block4_complete_3330_inst_req_0;
      WPIPE_Block4_complete_3330_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block4_complete_3330_inst_req_1;
      WPIPE_Block4_complete_3330_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_3332_wire_constant;
      Block4_complete_write_0_gI: SplitGuardInterface generic map(name => "Block4_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block4_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block4_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block4_complete_pipe_write_req(0),
          oack => Block4_complete_pipe_write_ack(0),
          odata => Block4_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_E_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_F is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block5_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block5_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block5_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block5_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block5_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block5_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_F;
architecture zeropad3D_F_arch of zeropad3D_F is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_F_CP_8333_start: Boolean;
  signal zeropad3D_F_CP_8333_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_3508_inst_ack_1 : boolean;
  signal phi_stmt_3503_req_1 : boolean;
  signal type_cast_3816_inst_req_0 : boolean;
  signal type_cast_3506_inst_ack_0 : boolean;
  signal type_cast_3752_inst_ack_0 : boolean;
  signal type_cast_3752_inst_req_0 : boolean;
  signal type_cast_3502_inst_req_1 : boolean;
  signal type_cast_3752_inst_req_1 : boolean;
  signal type_cast_3508_inst_req_1 : boolean;
  signal type_cast_3752_inst_ack_1 : boolean;
  signal if_stmt_3767_branch_req_0 : boolean;
  signal type_cast_3506_inst_req_0 : boolean;
  signal array_obj_ref_3740_index_offset_ack_1 : boolean;
  signal addr_of_3741_final_reg_ack_1 : boolean;
  signal array_obj_ref_3740_index_offset_req_1 : boolean;
  signal addr_of_3741_final_reg_req_1 : boolean;
  signal ptr_deref_3720_load_0_ack_1 : boolean;
  signal ptr_deref_3720_load_0_req_1 : boolean;
  signal type_cast_3508_inst_ack_0 : boolean;
  signal type_cast_3502_inst_ack_0 : boolean;
  signal type_cast_3508_inst_req_0 : boolean;
  signal phi_stmt_3503_ack_0 : boolean;
  signal array_obj_ref_3740_index_offset_ack_0 : boolean;
  signal phi_stmt_3497_req_0 : boolean;
  signal type_cast_3800_inst_ack_1 : boolean;
  signal type_cast_3816_inst_ack_0 : boolean;
  signal type_cast_3800_inst_req_1 : boolean;
  signal ptr_deref_3720_load_0_req_0 : boolean;
  signal type_cast_3502_inst_ack_1 : boolean;
  signal ptr_deref_3744_store_0_req_1 : boolean;
  signal type_cast_3842_inst_req_1 : boolean;
  signal type_cast_3842_inst_ack_1 : boolean;
  signal type_cast_3842_inst_ack_0 : boolean;
  signal phi_stmt_3497_req_1 : boolean;
  signal if_stmt_3767_branch_ack_1 : boolean;
  signal phi_stmt_3830_req_1 : boolean;
  signal ptr_deref_3744_store_0_ack_1 : boolean;
  signal type_cast_3816_inst_req_1 : boolean;
  signal type_cast_3734_inst_req_0 : boolean;
  signal type_cast_3816_inst_ack_1 : boolean;
  signal type_cast_3506_inst_req_1 : boolean;
  signal type_cast_3734_inst_ack_0 : boolean;
  signal type_cast_3842_inst_req_0 : boolean;
  signal if_stmt_3767_branch_ack_0 : boolean;
  signal type_cast_3506_inst_ack_1 : boolean;
  signal addr_of_3741_final_reg_req_0 : boolean;
  signal addr_of_3741_final_reg_ack_0 : boolean;
  signal phi_stmt_3837_req_1 : boolean;
  signal phi_stmt_3503_req_0 : boolean;
  signal RPIPE_Block5_starting_3341_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3341_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3341_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3341_inst_ack_1 : boolean;
  signal RPIPE_Block5_starting_3344_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3344_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3344_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3344_inst_ack_1 : boolean;
  signal RPIPE_Block5_starting_3347_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3347_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3347_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3347_inst_ack_1 : boolean;
  signal RPIPE_Block5_starting_3350_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3350_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3350_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3350_inst_ack_1 : boolean;
  signal RPIPE_Block5_starting_3353_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3353_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3353_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3353_inst_ack_1 : boolean;
  signal RPIPE_Block5_starting_3356_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3356_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3356_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3356_inst_ack_1 : boolean;
  signal RPIPE_Block5_starting_3359_inst_req_0 : boolean;
  signal RPIPE_Block5_starting_3359_inst_ack_0 : boolean;
  signal RPIPE_Block5_starting_3359_inst_req_1 : boolean;
  signal RPIPE_Block5_starting_3359_inst_ack_1 : boolean;
  signal type_cast_3364_inst_req_0 : boolean;
  signal type_cast_3364_inst_ack_0 : boolean;
  signal type_cast_3364_inst_req_1 : boolean;
  signal type_cast_3364_inst_ack_1 : boolean;
  signal type_cast_3374_inst_req_0 : boolean;
  signal type_cast_3374_inst_ack_0 : boolean;
  signal type_cast_3374_inst_req_1 : boolean;
  signal type_cast_3374_inst_ack_1 : boolean;
  signal type_cast_3384_inst_req_0 : boolean;
  signal type_cast_3384_inst_ack_0 : boolean;
  signal type_cast_3384_inst_req_1 : boolean;
  signal type_cast_3384_inst_ack_1 : boolean;
  signal type_cast_3388_inst_req_0 : boolean;
  signal type_cast_3388_inst_ack_0 : boolean;
  signal type_cast_3388_inst_req_1 : boolean;
  signal type_cast_3388_inst_ack_1 : boolean;
  signal type_cast_3392_inst_req_0 : boolean;
  signal type_cast_3392_inst_ack_0 : boolean;
  signal type_cast_3392_inst_req_1 : boolean;
  signal type_cast_3392_inst_ack_1 : boolean;
  signal type_cast_3396_inst_req_0 : boolean;
  signal type_cast_3396_inst_ack_0 : boolean;
  signal type_cast_3396_inst_req_1 : boolean;
  signal type_cast_3396_inst_ack_1 : boolean;
  signal type_cast_3405_inst_req_0 : boolean;
  signal type_cast_3405_inst_ack_0 : boolean;
  signal type_cast_3405_inst_req_1 : boolean;
  signal type_cast_3405_inst_ack_1 : boolean;
  signal type_cast_3409_inst_req_0 : boolean;
  signal type_cast_3409_inst_ack_0 : boolean;
  signal type_cast_3409_inst_req_1 : boolean;
  signal type_cast_3409_inst_ack_1 : boolean;
  signal type_cast_3439_inst_req_0 : boolean;
  signal type_cast_3439_inst_ack_0 : boolean;
  signal type_cast_3439_inst_req_1 : boolean;
  signal type_cast_3439_inst_ack_1 : boolean;
  signal type_cast_3513_inst_req_0 : boolean;
  signal type_cast_3513_inst_ack_0 : boolean;
  signal type_cast_3513_inst_req_1 : boolean;
  signal type_cast_3513_inst_ack_1 : boolean;
  signal if_stmt_3540_branch_req_0 : boolean;
  signal if_stmt_3540_branch_ack_1 : boolean;
  signal if_stmt_3540_branch_ack_0 : boolean;
  signal type_cast_3550_inst_req_0 : boolean;
  signal type_cast_3550_inst_ack_0 : boolean;
  signal type_cast_3550_inst_req_1 : boolean;
  signal type_cast_3550_inst_ack_1 : boolean;
  signal if_stmt_3577_branch_req_0 : boolean;
  signal ptr_deref_3720_load_0_ack_0 : boolean;
  signal array_obj_ref_3740_index_offset_req_0 : boolean;
  signal if_stmt_3577_branch_ack_1 : boolean;
  signal if_stmt_3577_branch_ack_0 : boolean;
  signal type_cast_3500_inst_ack_1 : boolean;
  signal type_cast_3800_inst_ack_0 : boolean;
  signal type_cast_3587_inst_req_0 : boolean;
  signal type_cast_3587_inst_ack_0 : boolean;
  signal type_cast_3800_inst_req_0 : boolean;
  signal type_cast_3587_inst_req_1 : boolean;
  signal type_cast_3587_inst_ack_1 : boolean;
  signal phi_stmt_3497_ack_0 : boolean;
  signal type_cast_3500_inst_req_1 : boolean;
  signal type_cast_3592_inst_req_0 : boolean;
  signal type_cast_3592_inst_ack_0 : boolean;
  signal type_cast_3592_inst_req_1 : boolean;
  signal type_cast_3592_inst_ack_1 : boolean;
  signal phi_stmt_3490_ack_0 : boolean;
  signal WPIPE_Block5_complete_3853_inst_ack_1 : boolean;
  signal WPIPE_Block5_complete_3853_inst_req_1 : boolean;
  signal type_cast_3626_inst_req_0 : boolean;
  signal type_cast_3626_inst_ack_0 : boolean;
  signal type_cast_3626_inst_req_1 : boolean;
  signal type_cast_3626_inst_ack_1 : boolean;
  signal phi_stmt_3490_req_1 : boolean;
  signal WPIPE_Block5_complete_3853_inst_ack_0 : boolean;
  signal WPIPE_Block5_complete_3853_inst_req_0 : boolean;
  signal ptr_deref_3744_store_0_ack_0 : boolean;
  signal ptr_deref_3744_store_0_req_0 : boolean;
  signal array_obj_ref_3632_index_offset_req_0 : boolean;
  signal array_obj_ref_3632_index_offset_ack_0 : boolean;
  signal array_obj_ref_3632_index_offset_req_1 : boolean;
  signal type_cast_3791_inst_ack_1 : boolean;
  signal array_obj_ref_3632_index_offset_ack_1 : boolean;
  signal type_cast_3500_inst_ack_0 : boolean;
  signal type_cast_3791_inst_req_1 : boolean;
  signal type_cast_3500_inst_req_0 : boolean;
  signal addr_of_3633_final_reg_req_0 : boolean;
  signal addr_of_3633_final_reg_ack_0 : boolean;
  signal addr_of_3633_final_reg_req_1 : boolean;
  signal type_cast_3791_inst_ack_0 : boolean;
  signal addr_of_3633_final_reg_ack_1 : boolean;
  signal type_cast_3496_inst_ack_1 : boolean;
  signal type_cast_3496_inst_req_1 : boolean;
  signal if_stmt_3823_branch_ack_0 : boolean;
  signal if_stmt_3823_branch_ack_1 : boolean;
  signal type_cast_3791_inst_req_0 : boolean;
  signal type_cast_3734_inst_ack_1 : boolean;
  signal type_cast_3734_inst_req_1 : boolean;
  signal ptr_deref_3636_store_0_req_0 : boolean;
  signal ptr_deref_3636_store_0_ack_0 : boolean;
  signal ptr_deref_3636_store_0_req_1 : boolean;
  signal ptr_deref_3636_store_0_ack_1 : boolean;
  signal type_cast_3496_inst_ack_0 : boolean;
  signal type_cast_3502_inst_req_0 : boolean;
  signal type_cast_3645_inst_req_0 : boolean;
  signal type_cast_3645_inst_ack_0 : boolean;
  signal phi_stmt_3490_req_0 : boolean;
  signal type_cast_3645_inst_req_1 : boolean;
  signal type_cast_3645_inst_ack_1 : boolean;
  signal if_stmt_3823_branch_req_0 : boolean;
  signal type_cast_3709_inst_req_0 : boolean;
  signal type_cast_3709_inst_ack_0 : boolean;
  signal type_cast_3709_inst_req_1 : boolean;
  signal type_cast_3709_inst_ack_1 : boolean;
  signal type_cast_3496_inst_req_0 : boolean;
  signal array_obj_ref_3715_index_offset_req_0 : boolean;
  signal array_obj_ref_3715_index_offset_ack_0 : boolean;
  signal array_obj_ref_3715_index_offset_req_1 : boolean;
  signal array_obj_ref_3715_index_offset_ack_1 : boolean;
  signal addr_of_3716_final_reg_req_0 : boolean;
  signal addr_of_3716_final_reg_ack_0 : boolean;
  signal addr_of_3716_final_reg_req_1 : boolean;
  signal addr_of_3716_final_reg_ack_1 : boolean;
  signal type_cast_3848_inst_req_0 : boolean;
  signal type_cast_3848_inst_ack_0 : boolean;
  signal type_cast_3848_inst_req_1 : boolean;
  signal type_cast_3848_inst_ack_1 : boolean;
  signal phi_stmt_3843_req_1 : boolean;
  signal type_cast_3833_inst_req_0 : boolean;
  signal type_cast_3833_inst_ack_0 : boolean;
  signal type_cast_3833_inst_req_1 : boolean;
  signal type_cast_3833_inst_ack_1 : boolean;
  signal phi_stmt_3830_req_0 : boolean;
  signal type_cast_3840_inst_req_0 : boolean;
  signal type_cast_3840_inst_ack_0 : boolean;
  signal type_cast_3840_inst_req_1 : boolean;
  signal type_cast_3840_inst_ack_1 : boolean;
  signal phi_stmt_3837_req_0 : boolean;
  signal type_cast_3846_inst_req_0 : boolean;
  signal type_cast_3846_inst_ack_0 : boolean;
  signal type_cast_3846_inst_req_1 : boolean;
  signal type_cast_3846_inst_ack_1 : boolean;
  signal phi_stmt_3843_req_0 : boolean;
  signal phi_stmt_3830_ack_0 : boolean;
  signal phi_stmt_3837_ack_0 : boolean;
  signal phi_stmt_3843_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_F_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_F_CP_8333_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_F_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_F_CP_8333_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_F_CP_8333_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_F_CP_8333_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_F_CP_8333: Block -- control-path 
    signal zeropad3D_F_CP_8333_elements: BooleanArray(138 downto 0);
    -- 
  begin -- 
    zeropad3D_F_CP_8333_elements(0) <= zeropad3D_F_CP_8333_start;
    zeropad3D_F_CP_8333_symbol <= zeropad3D_F_CP_8333_elements(90);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_3339/branch_block_stmt_3339__entry__
      -- CP-element group 0: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360__entry__
      -- CP-element group 0: 	 branch_block_stmt_3339/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/$entry
      -- CP-element group 0: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Sample/rr
      -- 
    rr_8399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(0), ack => RPIPE_Block5_starting_3341_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	138 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	100 
    -- CP-element group 1: 	102 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	105 
    -- CP-element group 1: 	106 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/merge_stmt_3829__exit__
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Sample/rr
      -- 
    cr_9269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(1), ack => type_cast_3508_inst_req_1); -- 
    rr_9264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(1), ack => type_cast_3508_inst_req_0); -- 
    cr_9292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(1), ack => type_cast_3500_inst_req_1); -- 
    rr_9287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(1), ack => type_cast_3500_inst_req_0); -- 
    cr_9315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(1), ack => type_cast_3496_inst_req_1); -- 
    rr_9310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(1), ack => type_cast_3496_inst_req_0); -- 
    zeropad3D_F_CP_8333_elements(1) <= zeropad3D_F_CP_8333_elements(138);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Update/cr
      -- 
    ra_8400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3341_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(2)); -- 
    cr_8404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(2), ack => RPIPE_Block5_starting_3341_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3341_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Sample/rr
      -- 
    ca_8405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3341_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(3)); -- 
    rr_8413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(3), ack => RPIPE_Block5_starting_3344_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_update_start_
      -- CP-element group 4: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Update/cr
      -- 
    ra_8414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3344_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(4)); -- 
    cr_8418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(4), ack => RPIPE_Block5_starting_3344_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3344_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Sample/rr
      -- 
    ca_8419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3344_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(5)); -- 
    rr_8427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(5), ack => RPIPE_Block5_starting_3347_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Update/cr
      -- 
    ra_8428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3347_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(6)); -- 
    cr_8432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(6), ack => RPIPE_Block5_starting_3347_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3347_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Sample/rr
      -- 
    ca_8433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3347_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(7)); -- 
    rr_8441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(7), ack => RPIPE_Block5_starting_3350_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_update_start_
      -- CP-element group 8: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Update/cr
      -- 
    ra_8442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3350_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(8)); -- 
    cr_8446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(8), ack => RPIPE_Block5_starting_3350_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3350_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Sample/rr
      -- 
    ca_8447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3350_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(9)); -- 
    rr_8455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(9), ack => RPIPE_Block5_starting_3353_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_update_start_
      -- CP-element group 10: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Update/cr
      -- 
    ra_8456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3353_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(10)); -- 
    cr_8460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(10), ack => RPIPE_Block5_starting_3353_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3353_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Sample/rr
      -- 
    ca_8461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3353_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(11)); -- 
    rr_8469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(11), ack => RPIPE_Block5_starting_3356_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_update_start_
      -- CP-element group 12: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Update/cr
      -- 
    ra_8470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3356_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(12)); -- 
    cr_8474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(12), ack => RPIPE_Block5_starting_3356_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3356_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Sample/rr
      -- 
    ca_8475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3356_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(13)); -- 
    rr_8483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(13), ack => RPIPE_Block5_starting_3359_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_update_start_
      -- CP-element group 14: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Update/cr
      -- 
    ra_8484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3359_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(14)); -- 
    cr_8488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(14), ack => RPIPE_Block5_starting_3359_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	32 
    -- CP-element group 15: 	33 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15:  members (61) 
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360__exit__
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487__entry__
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/$exit
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3342_to_assign_stmt_3360/RPIPE_Block5_starting_3359_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Update/cr
      -- 
    ca_8489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block5_starting_3359_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(15)); -- 
    rr_8500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3364_inst_req_0); -- 
    cr_8505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3364_inst_req_1); -- 
    rr_8514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3374_inst_req_0); -- 
    cr_8519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3374_inst_req_1); -- 
    rr_8528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3384_inst_req_0); -- 
    cr_8533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3384_inst_req_1); -- 
    rr_8542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3388_inst_req_0); -- 
    cr_8547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3388_inst_req_1); -- 
    rr_8556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3392_inst_req_0); -- 
    cr_8561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3392_inst_req_1); -- 
    rr_8570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3396_inst_req_0); -- 
    cr_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3396_inst_req_1); -- 
    rr_8584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3405_inst_req_0); -- 
    cr_8589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3405_inst_req_1); -- 
    rr_8598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3409_inst_req_0); -- 
    cr_8603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3409_inst_req_1); -- 
    rr_8612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3439_inst_req_0); -- 
    cr_8617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(15), ack => type_cast_3439_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Sample/ra
      -- 
    ra_8501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3364_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3364_Update/ca
      -- 
    ca_8506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3364_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Sample/ra
      -- 
    ra_8515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3374_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3374_Update/ca
      -- 
    ca_8520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3374_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Sample/ra
      -- 
    ra_8529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3384_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3384_Update/ca
      -- 
    ca_8534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3384_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Sample/ra
      -- 
    ra_8543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3388_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3388_Update/ca
      -- 
    ca_8548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3388_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Sample/ra
      -- 
    ra_8557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3392_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3392_Update/ca
      -- 
    ca_8562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3392_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Sample/ra
      -- 
    ra_8571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3396_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3396_Update/ca
      -- 
    ca_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3396_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Sample/ra
      -- 
    ra_8585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3405_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3405_Update/ca
      -- 
    ca_8590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3405_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Sample/ra
      -- 
    ra_8599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3409_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3409_Update/ca
      -- 
    ca_8604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3409_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Sample/ra
      -- 
    ra_8613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3439_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/type_cast_3439_Update/ca
      -- 
    ca_8618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3439_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	91 
    -- CP-element group 34: 	92 
    -- CP-element group 34: 	94 
    -- CP-element group 34: 	95 
    -- CP-element group 34: 	97 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487__exit__
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3490/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/assign_stmt_3365_to_assign_stmt_3487/$exit
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/$entry
      -- CP-element group 34: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/$entry
      -- 
    cr_9235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(34), ack => type_cast_3502_inst_req_1); -- 
    rr_9207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(34), ack => type_cast_3506_inst_req_0); -- 
    cr_9212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(34), ack => type_cast_3506_inst_req_1); -- 
    rr_9230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(34), ack => type_cast_3502_inst_req_0); -- 
    zeropad3D_F_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(29) & zeropad3D_F_CP_8333_elements(31) & zeropad3D_F_CP_8333_elements(33) & zeropad3D_F_CP_8333_elements(23) & zeropad3D_F_CP_8333_elements(21) & zeropad3D_F_CP_8333_elements(25) & zeropad3D_F_CP_8333_elements(27) & zeropad3D_F_CP_8333_elements(17) & zeropad3D_F_CP_8333_elements(19);
      gj_zeropad3D_F_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	113 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Sample/ra
      -- 
    ra_8630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3513_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	113 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (13) 
      -- CP-element group 36: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539__exit__
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540__entry__
      -- CP-element group 36: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/$exit
      -- CP-element group 36: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_3339/R_orx_xcond_3541_place
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_3339/if_stmt_3540_else_link/$entry
      -- 
    ca_8635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3513_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(36)); -- 
    branch_req_8643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(36), ack => if_stmt_3540_branch_req_0); -- 
    -- CP-element group 37:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	40 
    -- CP-element group 37:  members (18) 
      -- CP-element group 37: 	 branch_block_stmt_3339/merge_stmt_3546_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_3339/merge_stmt_3546_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_3339/whilex_xbody_lorx_xlhsx_xfalse65_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_3339/whilex_xbody_lorx_xlhsx_xfalse65_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_3339/merge_stmt_3546__exit__
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576__entry__
      -- CP-element group 37: 	 branch_block_stmt_3339/merge_stmt_3546_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_3339/merge_stmt_3546_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_3339/if_stmt_3540_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_3339/if_stmt_3540_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_3339/whilex_xbody_lorx_xlhsx_xfalse65
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/$entry
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_update_start_
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Update/cr
      -- 
    if_choice_transition_8648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3540_branch_ack_1, ack => zeropad3D_F_CP_8333_elements(37)); -- 
    rr_8665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(37), ack => type_cast_3550_inst_req_0); -- 
    cr_8670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(37), ack => type_cast_3550_inst_req_1); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	114 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_3339/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 38: 	 branch_block_stmt_3339/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_3339/if_stmt_3540_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_3339/if_stmt_3540_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_3339/whilex_xbody_ifx_xthen
      -- 
    else_choice_transition_8652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3540_branch_ack_0, ack => zeropad3D_F_CP_8333_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Sample/ra
      -- 
    ra_8666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3550_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(39)); -- 
    -- CP-element group 40:  branch  transition  place  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (13) 
      -- CP-element group 40: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576__exit__
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577__entry__
      -- CP-element group 40: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/$exit
      -- CP-element group 40: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_3339/assign_stmt_3551_to_assign_stmt_3576/type_cast_3550_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577_dead_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577_eval_test/$entry
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577_eval_test/$exit
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577_eval_test/branch_req
      -- CP-element group 40: 	 branch_block_stmt_3339/R_orx_xcond196_3578_place
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577_if_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_3339/if_stmt_3577_else_link/$entry
      -- 
    ca_8671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3550_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(40)); -- 
    branch_req_8679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(40), ack => if_stmt_3577_branch_req_0); -- 
    -- CP-element group 41:  fork  transition  place  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	58 
    -- CP-element group 41: 	60 
    -- CP-element group 41: 	62 
    -- CP-element group 41: 	64 
    -- CP-element group 41: 	66 
    -- CP-element group 41: 	68 
    -- CP-element group 41: 	70 
    -- CP-element group 41: 	72 
    -- CP-element group 41: 	75 
    -- CP-element group 41:  members (46) 
      -- CP-element group 41: 	 branch_block_stmt_3339/merge_stmt_3641_PhiReqMerge
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_complete/req
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/merge_stmt_3641_PhiAck/dummy
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746__entry__
      -- CP-element group 41: 	 branch_block_stmt_3339/merge_stmt_3641__exit__
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_3339/lorx_xlhsx_xfalse65_ifx_xelse_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/lorx_xlhsx_xfalse65_ifx_xelse_PhiReq/$exit
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/merge_stmt_3641_PhiAck/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/merge_stmt_3641_PhiAck/$exit
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/if_stmt_3577_if_link/$exit
      -- CP-element group 41: 	 branch_block_stmt_3339/if_stmt_3577_if_link/if_choice_transition
      -- CP-element group 41: 	 branch_block_stmt_3339/lorx_xlhsx_xfalse65_ifx_xelse
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_complete/req
      -- CP-element group 41: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_update_start_
      -- 
    if_choice_transition_8684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3577_branch_ack_1, ack => zeropad3D_F_CP_8333_elements(41)); -- 
    req_9002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => array_obj_ref_3740_index_offset_req_1); -- 
    req_9017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => addr_of_3741_final_reg_req_1); -- 
    cr_8952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => ptr_deref_3720_load_0_req_1); -- 
    cr_9067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => ptr_deref_3744_store_0_req_1); -- 
    cr_8971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => type_cast_3734_inst_req_1); -- 
    rr_8842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => type_cast_3645_inst_req_0); -- 
    cr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => type_cast_3645_inst_req_1); -- 
    cr_8861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => type_cast_3709_inst_req_1); -- 
    req_8892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => array_obj_ref_3715_index_offset_req_1); -- 
    req_8907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(41), ack => addr_of_3716_final_reg_req_1); -- 
    -- CP-element group 42:  transition  place  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	114 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_3339/lorx_xlhsx_xfalse65_ifx_xthen_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_3339/lorx_xlhsx_xfalse65_ifx_xthen_PhiReq/$exit
      -- CP-element group 42: 	 branch_block_stmt_3339/if_stmt_3577_else_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_3339/if_stmt_3577_else_link/else_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_3339/lorx_xlhsx_xfalse65_ifx_xthen
      -- 
    else_choice_transition_8688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3577_branch_ack_0, ack => zeropad3D_F_CP_8333_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	114 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Sample/ra
      -- 
    ra_8702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3587_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	114 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Update/ca
      -- 
    ca_8707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3587_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	114 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Sample/ra
      -- 
    ra_8716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3592_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	114 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Update/ca
      -- 
    ca_8721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3592_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Sample/rr
      -- 
    rr_8729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(47), ack => type_cast_3626_inst_req_0); -- 
    zeropad3D_F_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(44) & zeropad3D_F_CP_8333_elements(46);
      gj_zeropad3D_F_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Sample/ra
      -- 
    ra_8730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3626_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	114 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Sample/req
      -- 
    ca_8735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3626_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(49)); -- 
    req_8760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(49), ack => array_obj_ref_3632_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	56 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Sample/ack
      -- 
    ack_8761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3632_index_offset_ack_0, ack => zeropad3D_F_CP_8333_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	114 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_request/req
      -- 
    ack_8766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3632_index_offset_ack_1, ack => zeropad3D_F_CP_8333_elements(51)); -- 
    req_8775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(51), ack => addr_of_3633_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_request/ack
      -- 
    ack_8776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3633_final_reg_ack_0, ack => zeropad3D_F_CP_8333_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	114 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (28) 
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/ptr_deref_3636_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/ptr_deref_3636_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/ptr_deref_3636_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/ptr_deref_3636_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/word_access_start/word_0/rr
      -- 
    ack_8781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3633_final_reg_ack_1, ack => zeropad3D_F_CP_8333_elements(53)); -- 
    rr_8819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(53), ack => ptr_deref_3636_store_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Sample/word_access_start/word_0/ra
      -- 
    ra_8820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3636_store_0_ack_0, ack => zeropad3D_F_CP_8333_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	114 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/word_access_complete/word_0/ca
      -- 
    ca_8831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3636_store_0_ack_1, ack => zeropad3D_F_CP_8333_elements(55)); -- 
    -- CP-element group 56:  join  transition  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	50 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	115 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639__exit__
      -- CP-element group 56: 	 branch_block_stmt_3339/ifx_xthen_ifx_xend
      -- CP-element group 56: 	 branch_block_stmt_3339/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_3339/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/$exit
      -- 
    zeropad3D_F_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(55) & zeropad3D_F_CP_8333_elements(50);
      gj_zeropad3D_F_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Sample/ra
      -- 
    ra_8843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3645_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	67 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3645_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Sample/rr
      -- 
    ca_8848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3645_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(58)); -- 
    rr_8856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(58), ack => type_cast_3709_inst_req_0); -- 
    rr_8966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(58), ack => type_cast_3734_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Sample/ra
      -- 
    ra_8857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3709_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	41 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (16) 
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3709_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_scale_1/scale_rename_req
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Sample/req
      -- 
    ca_8862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3709_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(60)); -- 
    req_8887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(60), ack => array_obj_ref_3715_index_offset_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	76 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Sample/ack
      -- 
    ack_8888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3715_index_offset_ack_0, ack => zeropad3D_F_CP_8333_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	41 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (11) 
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_offset_calculated
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_final_index_sum_regn_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3715_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_request/$entry
      -- CP-element group 62: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_request/req
      -- 
    ack_8893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3715_index_offset_ack_1, ack => zeropad3D_F_CP_8333_elements(62)); -- 
    req_8902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(62), ack => addr_of_3716_final_reg_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_request/$exit
      -- CP-element group 63: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_request/ack
      -- 
    ack_8903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3716_final_reg_ack_0, ack => zeropad3D_F_CP_8333_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	41 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (24) 
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/word_access_start/word_0/rr
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3716_complete/ack
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_word_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_address_resized
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_addr_resize/$entry
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_addr_resize/$exit
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_addr_resize/base_resize_req
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_addr_resize/base_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_word_addrgen/$entry
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_word_addrgen/$exit
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_word_addrgen/root_register_req
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_word_addrgen/root_register_ack
      -- CP-element group 64: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/$entry
      -- 
    ack_8908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3716_final_reg_ack_1, ack => zeropad3D_F_CP_8333_elements(64)); -- 
    rr_8941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(64), ack => ptr_deref_3720_load_0_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/word_access_start/word_0/ra
      -- CP-element group 65: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Sample/$exit
      -- 
    ra_8942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3720_load_0_ack_0, ack => zeropad3D_F_CP_8333_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	41 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	73 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/ptr_deref_3720_Merge/$exit
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/ptr_deref_3720_Merge/$entry
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/word_access_complete/word_0/ca
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/ptr_deref_3720_Merge/merge_ack
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/ptr_deref_3720_Merge/merge_req
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3720_update_completed_
      -- 
    ca_8953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3720_load_0_ack_1, ack => zeropad3D_F_CP_8333_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	58 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Sample/ra
      -- 
    ra_8967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3734_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	41 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_scaled_1
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_resized_1
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_computed_1
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_scale_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_resize_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_resize_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_resize_1/index_resize_req
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_resize_1/index_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_scale_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Sample/req
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/type_cast_3734_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_scale_1/scale_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_index_scale_1/scale_rename_req
      -- 
    ca_8972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3734_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(68)); -- 
    req_8997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(68), ack => array_obj_ref_3740_index_offset_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	76 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_sample_complete
      -- 
    ack_8998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3740_index_offset_ack_0, ack => zeropad3D_F_CP_8333_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	41 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (11) 
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_offset_calculated
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_final_index_sum_regn_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_request/$entry
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_request/req
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/array_obj_ref_3740_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_sample_start_
      -- 
    ack_9003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3740_index_offset_ack_1, ack => zeropad3D_F_CP_8333_elements(70)); -- 
    req_9012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(70), ack => addr_of_3741_final_reg_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_request/$exit
      -- CP-element group 71: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_request/ack
      -- CP-element group 71: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_sample_completed_
      -- 
    ack_9013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3741_final_reg_ack_0, ack => zeropad3D_F_CP_8333_elements(71)); -- 
    -- CP-element group 72:  fork  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	41 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (19) 
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_complete/ack
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/addr_of_3741_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_word_addrgen/root_register_ack
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_word_address_calculated
      -- 
    ack_9018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3741_final_reg_ack_1, ack => zeropad3D_F_CP_8333_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/ptr_deref_3744_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/ptr_deref_3744_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/ptr_deref_3744_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/ptr_deref_3744_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/$entry
      -- 
    rr_9056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(73), ack => ptr_deref_3744_store_0_req_0); -- 
    zeropad3D_F_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(66) & zeropad3D_F_CP_8333_elements(72);
      gj_zeropad3D_F_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/word_access_start/word_0/ra
      -- CP-element group 74: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Sample/$exit
      -- 
    ra_9057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3744_store_0_ack_0, ack => zeropad3D_F_CP_8333_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_Update/word_access_complete/word_0/ca
      -- CP-element group 75: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/ptr_deref_3744_update_completed_
      -- 
    ca_9068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3744_store_0_ack_1, ack => zeropad3D_F_CP_8333_elements(75)); -- 
    -- CP-element group 76:  join  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	61 
    -- CP-element group 76: 	69 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	115 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746__exit__
      -- CP-element group 76: 	 branch_block_stmt_3339/ifx_xelse_ifx_xend
      -- CP-element group 76: 	 branch_block_stmt_3339/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_3339/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_3339/assign_stmt_3646_to_assign_stmt_3746/$exit
      -- 
    zeropad3D_F_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(61) & zeropad3D_F_CP_8333_elements(69) & zeropad3D_F_CP_8333_elements(75);
      gj_zeropad3D_F_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	115 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_sample_completed_
      -- 
    ra_9080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3752_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(77)); -- 
    -- CP-element group 78:  branch  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	115 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (13) 
      -- CP-element group 78: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767_eval_test/branch_req
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767_dead_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767_eval_test/$exit
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767_eval_test/$entry
      -- CP-element group 78: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767_if_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767__entry__
      -- CP-element group 78: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766__exit__
      -- CP-element group 78: 	 branch_block_stmt_3339/if_stmt_3767_else_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/$exit
      -- CP-element group 78: 	 branch_block_stmt_3339/R_cmp149_3768_place
      -- 
    ca_9085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3752_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(78)); -- 
    branch_req_9093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(78), ack => if_stmt_3767_branch_req_0); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	124 
    -- CP-element group 79: 	125 
    -- CP-element group 79: 	127 
    -- CP-element group 79: 	128 
    -- CP-element group 79: 	130 
    -- CP-element group 79: 	131 
    -- CP-element group 79:  members (40) 
      -- CP-element group 79: 	 branch_block_stmt_3339/assign_stmt_3779__entry__
      -- CP-element group 79: 	 branch_block_stmt_3339/merge_stmt_3773__exit__
      -- CP-element group 79: 	 branch_block_stmt_3339/assign_stmt_3779__exit__
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190
      -- CP-element group 79: 	 branch_block_stmt_3339/if_stmt_3767_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xend_ifx_xthen151_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xend_ifx_xthen151_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_3339/if_stmt_3767_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_3339/merge_stmt_3773_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_3339/merge_stmt_3773_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/merge_stmt_3773_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_3339/merge_stmt_3773_PhiAck/dummy
      -- CP-element group 79: 	 branch_block_stmt_3339/assign_stmt_3779/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/assign_stmt_3779/$exit
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xend_ifx_xthen151
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Update/cr
      -- 
    if_choice_transition_9098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3767_branch_ack_1, ack => zeropad3D_F_CP_8333_elements(79)); -- 
    rr_9470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(79), ack => type_cast_3833_inst_req_0); -- 
    cr_9475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(79), ack => type_cast_3833_inst_req_1); -- 
    rr_9493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(79), ack => type_cast_3840_inst_req_0); -- 
    cr_9498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(79), ack => type_cast_3840_inst_req_1); -- 
    rr_9516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(79), ack => type_cast_3846_inst_req_0); -- 
    cr_9521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(79), ack => type_cast_3846_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  place  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80: 	84 
    -- CP-element group 80: 	86 
    -- CP-element group 80:  members (24) 
      -- CP-element group 80: 	 branch_block_stmt_3339/ifx_xend_ifx_xelse156
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_update_start_
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_3339/merge_stmt_3781__exit__
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822__entry__
      -- CP-element group 80: 	 branch_block_stmt_3339/if_stmt_3767_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_3339/merge_stmt_3781_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_3339/ifx_xend_ifx_xelse156_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_3339/ifx_xend_ifx_xelse156_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_3339/if_stmt_3767_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_3339/merge_stmt_3781_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_3339/merge_stmt_3781_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_3339/merge_stmt_3781_PhiAck/dummy
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_update_start_
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_update_start_
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/$entry
      -- 
    else_choice_transition_9102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3767_branch_ack_0, ack => zeropad3D_F_CP_8333_elements(80)); -- 
    cr_9137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(80), ack => type_cast_3800_inst_req_1); -- 
    cr_9151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(80), ack => type_cast_3816_inst_req_1); -- 
    cr_9123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(80), ack => type_cast_3791_inst_req_1); -- 
    rr_9118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(80), ack => type_cast_3791_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_sample_completed_
      -- 
    ra_9119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3791_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3791_update_completed_
      -- 
    ca_9124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3791_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(82)); -- 
    rr_9132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(82), ack => type_cast_3800_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_sample_completed_
      -- 
    ra_9133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3800_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3800_update_completed_
      -- 
    ca_9138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3800_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(84)); -- 
    rr_9146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(84), ack => type_cast_3816_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Sample/ra
      -- 
    ra_9147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3816_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(85)); -- 
    -- CP-element group 86:  branch  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	80 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (13) 
      -- CP-element group 86: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_3339/R_cmp182_3824_place
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823__entry__
      -- CP-element group 86: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822__exit__
      -- CP-element group 86: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/type_cast_3816_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823_else_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_3339/assign_stmt_3787_to_assign_stmt_3822/$exit
      -- CP-element group 86: 	 branch_block_stmt_3339/if_stmt_3823_eval_test/$entry
      -- 
    ca_9152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3816_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(86)); -- 
    branch_req_9160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(86), ack => if_stmt_3823_branch_req_0); -- 
    -- CP-element group 87:  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (15) 
      -- CP-element group 87: 	 branch_block_stmt_3339/ifx_xelse156_whilex_xend
      -- CP-element group 87: 	 branch_block_stmt_3339/merge_stmt_3851_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_3339/merge_stmt_3851__exit__
      -- CP-element group 87: 	 branch_block_stmt_3339/assign_stmt_3856__entry__
      -- CP-element group 87: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_3339/assign_stmt_3856/$entry
      -- CP-element group 87: 	 branch_block_stmt_3339/if_stmt_3823_if_link/if_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_3339/if_stmt_3823_if_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_3339/ifx_xelse156_whilex_xend_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_3339/ifx_xelse156_whilex_xend_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_3339/merge_stmt_3851_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_3339/merge_stmt_3851_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_3339/merge_stmt_3851_PhiAck/dummy
      -- 
    if_choice_transition_9165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3823_branch_ack_1, ack => zeropad3D_F_CP_8333_elements(87)); -- 
    req_9182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(87), ack => WPIPE_Block5_complete_3853_inst_req_0); -- 
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	116 
    -- CP-element group 88: 	117 
    -- CP-element group 88: 	118 
    -- CP-element group 88: 	120 
    -- CP-element group 88: 	121 
    -- CP-element group 88:  members (22) 
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3830/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/if_stmt_3823_else_link/else_choice_transition
      -- CP-element group 88: 	 branch_block_stmt_3339/if_stmt_3823_else_link/$exit
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Update/cr
      -- 
    else_choice_transition_9169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3823_branch_ack_0, ack => zeropad3D_F_CP_8333_elements(88)); -- 
    cr_9426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(88), ack => type_cast_3842_inst_req_1); -- 
    rr_9421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(88), ack => type_cast_3842_inst_req_0); -- 
    rr_9444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(88), ack => type_cast_3848_inst_req_0); -- 
    cr_9449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(88), ack => type_cast_3848_inst_req_1); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Update/req
      -- CP-element group 89: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_update_start_
      -- CP-element group 89: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_sample_completed_
      -- 
    ack_9183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_complete_3853_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(89)); -- 
    req_9187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(89), ack => WPIPE_Block5_complete_3853_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (16) 
      -- CP-element group 90: 	 branch_block_stmt_3339/$exit
      -- CP-element group 90: 	 branch_block_stmt_3339/branch_block_stmt_3339__exit__
      -- CP-element group 90: 	 $exit
      -- CP-element group 90: 	 branch_block_stmt_3339/merge_stmt_3858_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_3339/assign_stmt_3856__exit__
      -- CP-element group 90: 	 branch_block_stmt_3339/return__
      -- CP-element group 90: 	 branch_block_stmt_3339/merge_stmt_3858__exit__
      -- CP-element group 90: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_3339/assign_stmt_3856/WPIPE_Block5_complete_3853_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_3339/assign_stmt_3856/$exit
      -- CP-element group 90: 	 branch_block_stmt_3339/return___PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_3339/return___PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_3339/merge_stmt_3858_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_3339/merge_stmt_3858_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_3339/merge_stmt_3858_PhiAck/dummy
      -- 
    ack_9188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block5_complete_3853_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	34 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Sample/ra
      -- 
    ra_9208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3506_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	34 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/Update/ca
      -- 
    ca_9213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3506_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	98 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/$exit
      -- CP-element group 93: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/$exit
      -- CP-element group 93: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3506/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_req
      -- 
    phi_stmt_3503_req_9214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3503_req_9214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(93), ack => phi_stmt_3503_req_0); -- 
    zeropad3D_F_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(91) & zeropad3D_F_CP_8333_elements(92);
      gj_zeropad3D_F_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	34 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Sample/$exit
      -- 
    ra_9231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3502_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	34 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/Update/ca
      -- 
    ca_9236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3502_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/$exit
      -- CP-element group 96: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/$exit
      -- CP-element group 96: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_req
      -- CP-element group 96: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3502/SplitProtocol/$exit
      -- 
    phi_stmt_3497_req_9237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3497_req_9237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(96), ack => phi_stmt_3497_req_1); -- 
    zeropad3D_F_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(94) & zeropad3D_F_CP_8333_elements(95);
      gj_zeropad3D_F_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  output  delay-element  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	34 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3490/$exit
      -- CP-element group 97: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_req
      -- CP-element group 97: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3494_konst_delay_trans
      -- CP-element group 97: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/$exit
      -- 
    phi_stmt_3490_req_9245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3490_req_9245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(97), ack => phi_stmt_3490_req_0); -- 
    -- Element group zeropad3D_F_CP_8333_elements(97) is a control-delay.
    cp_element_97_delay: control_delay_element  generic map(name => " 97_delay", delay_value => 1)  port map(req => zeropad3D_F_CP_8333_elements(34), ack => zeropad3D_F_CP_8333_elements(97), clk => clk, reset =>reset);
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	93 
    -- CP-element group 98: 	96 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	109 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_3339/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_F_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_F_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(93) & zeropad3D_F_CP_8333_elements(96) & zeropad3D_F_CP_8333_elements(97);
      gj_zeropad3D_F_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Sample/$exit
      -- 
    ra_9265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3508_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Update/ca
      -- CP-element group 100: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/Update/$exit
      -- 
    ca_9270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3508_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_req
      -- CP-element group 101: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/type_cast_3508/$exit
      -- CP-element group 101: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/phi_stmt_3503_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3503/$exit
      -- 
    phi_stmt_3503_req_9271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3503_req_9271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(101), ack => phi_stmt_3503_req_1); -- 
    zeropad3D_F_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(99) & zeropad3D_F_CP_8333_elements(100);
      gj_zeropad3D_F_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Sample/$exit
      -- 
    ra_9288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3500_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Update/ca
      -- CP-element group 103: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/Update/$exit
      -- 
    ca_9293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3500_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/$exit
      -- CP-element group 104: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_req
      -- CP-element group 104: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/$exit
      -- CP-element group 104: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3497/phi_stmt_3497_sources/type_cast_3500/SplitProtocol/$exit
      -- 
    phi_stmt_3497_req_9294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3497_req_9294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(104), ack => phi_stmt_3497_req_0); -- 
    zeropad3D_F_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(102) & zeropad3D_F_CP_8333_elements(103);
      gj_zeropad3D_F_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	1 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Sample/ra
      -- 
    ra_9311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3496_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/Update/$exit
      -- 
    ca_9316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3496_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/$exit
      -- CP-element group 107: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/$exit
      -- CP-element group 107: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_sources/type_cast_3496/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/phi_stmt_3490/phi_stmt_3490_req
      -- 
    phi_stmt_3490_req_9317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3490_req_9317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(107), ack => phi_stmt_3490_req_1); -- 
    zeropad3D_F_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(105) & zeropad3D_F_CP_8333_elements(106);
      gj_zeropad3D_F_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_3339/ifx_xend190_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_F_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(101) & zeropad3D_F_CP_8333_elements(104) & zeropad3D_F_CP_8333_elements(107);
      gj_zeropad3D_F_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	98 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_3339/merge_stmt_3489_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_3339/merge_stmt_3489_PhiAck/$entry
      -- 
    zeropad3D_F_CP_8333_elements(109) <= OrReduce(zeropad3D_F_CP_8333_elements(98) & zeropad3D_F_CP_8333_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_3339/merge_stmt_3489_PhiAck/phi_stmt_3490_ack
      -- 
    phi_stmt_3490_ack_9322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3490_ack_0, ack => zeropad3D_F_CP_8333_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_3339/merge_stmt_3489_PhiAck/phi_stmt_3497_ack
      -- 
    phi_stmt_3497_ack_9323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3497_ack_0, ack => zeropad3D_F_CP_8333_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_3339/merge_stmt_3489_PhiAck/phi_stmt_3503_ack
      -- 
    phi_stmt_3503_ack_9324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3503_ack_0, ack => zeropad3D_F_CP_8333_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	35 
    -- CP-element group 113: 	36 
    -- CP-element group 113:  members (10) 
      -- CP-element group 113: 	 branch_block_stmt_3339/merge_stmt_3489__exit__
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539__entry__
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/$entry
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_update_start_
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_3339/assign_stmt_3514_to_assign_stmt_3539/type_cast_3513_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_3339/merge_stmt_3489_PhiAck/$exit
      -- 
    rr_8629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(113), ack => type_cast_3513_inst_req_0); -- 
    cr_8634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(113), ack => type_cast_3513_inst_req_1); -- 
    zeropad3D_F_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(110) & zeropad3D_F_CP_8333_elements(111) & zeropad3D_F_CP_8333_elements(112);
      gj_zeropad3D_F_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  merge  fork  transition  place  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	38 
    -- CP-element group 114: 	42 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	55 
    -- CP-element group 114: 	43 
    -- CP-element group 114: 	44 
    -- CP-element group 114: 	45 
    -- CP-element group 114: 	46 
    -- CP-element group 114: 	49 
    -- CP-element group 114: 	51 
    -- CP-element group 114: 	53 
    -- CP-element group 114:  members (33) 
      -- CP-element group 114: 	 branch_block_stmt_3339/merge_stmt_3583_PhiReqMerge
      -- CP-element group 114: 	 branch_block_stmt_3339/merge_stmt_3583__exit__
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639__entry__
      -- CP-element group 114: 	 branch_block_stmt_3339/merge_stmt_3583_PhiAck/dummy
      -- CP-element group 114: 	 branch_block_stmt_3339/merge_stmt_3583_PhiAck/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/merge_stmt_3583_PhiAck/$exit
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_update_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3587_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_update_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3592_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_update_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/type_cast_3626_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_update_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_update_start
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/array_obj_ref_3632_final_index_sum_regn_Update/req
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/addr_of_3633_complete/req
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_update_start_
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/word_access_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/word_access_complete/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_3339/assign_stmt_3588_to_assign_stmt_3639/ptr_deref_3636_Update/word_access_complete/word_0/cr
      -- 
    rr_8701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => type_cast_3587_inst_req_0); -- 
    cr_8706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => type_cast_3587_inst_req_1); -- 
    rr_8715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => type_cast_3592_inst_req_0); -- 
    cr_8720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => type_cast_3592_inst_req_1); -- 
    cr_8734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => type_cast_3626_inst_req_1); -- 
    req_8765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => array_obj_ref_3632_index_offset_req_1); -- 
    req_8780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => addr_of_3633_final_reg_req_1); -- 
    cr_8830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(114), ack => ptr_deref_3636_store_0_req_1); -- 
    zeropad3D_F_CP_8333_elements(114) <= OrReduce(zeropad3D_F_CP_8333_elements(38) & zeropad3D_F_CP_8333_elements(42));
    -- CP-element group 115:  merge  fork  transition  place  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	56 
    -- CP-element group 115: 	76 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	77 
    -- CP-element group 115: 	78 
    -- CP-element group 115:  members (13) 
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_3339/merge_stmt_3748__exit__
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766__entry__
      -- CP-element group 115: 	 branch_block_stmt_3339/merge_stmt_3748_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_3339/merge_stmt_3748_PhiAck/dummy
      -- CP-element group 115: 	 branch_block_stmt_3339/merge_stmt_3748_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_3339/merge_stmt_3748_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_update_start_
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/type_cast_3752_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_3339/assign_stmt_3753_to_assign_stmt_3766/$entry
      -- 
    rr_9079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(115), ack => type_cast_3752_inst_req_0); -- 
    cr_9084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(115), ack => type_cast_3752_inst_req_1); -- 
    zeropad3D_F_CP_8333_elements(115) <= OrReduce(zeropad3D_F_CP_8333_elements(56) & zeropad3D_F_CP_8333_elements(76));
    -- CP-element group 116:  transition  output  delay-element  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	88 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	123 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3830/$exit
      -- CP-element group 116: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_req
      -- CP-element group 116: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3836_konst_delay_trans
      -- 
    phi_stmt_3830_req_9405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3830_req_9405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(116), ack => phi_stmt_3830_req_1); -- 
    -- Element group zeropad3D_F_CP_8333_elements(116) is a control-delay.
    cp_element_116_delay: control_delay_element  generic map(name => " 116_delay", delay_value => 1)  port map(req => zeropad3D_F_CP_8333_elements(88), ack => zeropad3D_F_CP_8333_elements(116), clk => clk, reset =>reset);
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	88 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Sample/$exit
      -- 
    ra_9422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3842_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Update/ca
      -- CP-element group 118: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/Update/$exit
      -- 
    ca_9427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3842_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/$exit
      -- CP-element group 119: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_req
      -- CP-element group 119: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3842/$exit
      -- CP-element group 119: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/$exit
      -- 
    phi_stmt_3837_req_9428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3837_req_9428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(119), ack => phi_stmt_3837_req_1); -- 
    zeropad3D_F_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(117) & zeropad3D_F_CP_8333_elements(118);
      gj_zeropad3D_F_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	88 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Sample/ra
      -- 
    ra_9445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3848_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	88 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/Update/ca
      -- 
    ca_9450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3848_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/$exit
      -- CP-element group 122: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/$exit
      -- CP-element group 122: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3848/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_req
      -- 
    phi_stmt_3843_req_9451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3843_req_9451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(122), ack => phi_stmt_3843_req_1); -- 
    zeropad3D_F_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(120) & zeropad3D_F_CP_8333_elements(121);
      gj_zeropad3D_F_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	116 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	134 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_3339/ifx_xelse156_ifx_xend190_PhiReq/$exit
      -- 
    zeropad3D_F_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(116) & zeropad3D_F_CP_8333_elements(119) & zeropad3D_F_CP_8333_elements(122);
      gj_zeropad3D_F_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	79 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Sample/ra
      -- 
    ra_9471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3833_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/Update/ca
      -- 
    ca_9476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3833_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	133 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/$exit
      -- CP-element group 126: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/$exit
      -- CP-element group 126: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_sources/type_cast_3833/SplitProtocol/$exit
      -- CP-element group 126: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3830/phi_stmt_3830_req
      -- 
    phi_stmt_3830_req_9477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3830_req_9477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(126), ack => phi_stmt_3830_req_0); -- 
    zeropad3D_F_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(124) & zeropad3D_F_CP_8333_elements(125);
      gj_zeropad3D_F_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	79 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Sample/ra
      -- 
    ra_9494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3840_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	79 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/Update/ca
      -- 
    ca_9499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3840_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/$exit
      -- CP-element group 129: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/$exit
      -- CP-element group 129: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/$exit
      -- CP-element group 129: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_sources/type_cast_3840/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3837/phi_stmt_3837_req
      -- 
    phi_stmt_3837_req_9500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3837_req_9500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(129), ack => phi_stmt_3837_req_0); -- 
    zeropad3D_F_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(127) & zeropad3D_F_CP_8333_elements(128);
      gj_zeropad3D_F_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	79 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Sample/ra
      -- 
    ra_9517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3846_inst_ack_0, ack => zeropad3D_F_CP_8333_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	79 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/Update/ca
      -- 
    ca_9522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3846_inst_ack_1, ack => zeropad3D_F_CP_8333_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/$exit
      -- CP-element group 132: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/$exit
      -- CP-element group 132: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/$exit
      -- CP-element group 132: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_sources/type_cast_3846/SplitProtocol/$exit
      -- CP-element group 132: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/phi_stmt_3843/phi_stmt_3843_req
      -- 
    phi_stmt_3843_req_9523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3843_req_9523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_F_CP_8333_elements(132), ack => phi_stmt_3843_req_0); -- 
    zeropad3D_F_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(130) & zeropad3D_F_CP_8333_elements(131);
      gj_zeropad3D_F_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	126 
    -- CP-element group 133: 	129 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_3339/ifx_xthen151_ifx_xend190_PhiReq/$exit
      -- 
    zeropad3D_F_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(126) & zeropad3D_F_CP_8333_elements(129) & zeropad3D_F_CP_8333_elements(132);
      gj_zeropad3D_F_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  merge  fork  transition  place  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	123 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_3339/merge_stmt_3829_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_3339/merge_stmt_3829_PhiAck/$entry
      -- 
    zeropad3D_F_CP_8333_elements(134) <= OrReduce(zeropad3D_F_CP_8333_elements(123) & zeropad3D_F_CP_8333_elements(133));
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_3339/merge_stmt_3829_PhiAck/phi_stmt_3830_ack
      -- 
    phi_stmt_3830_ack_9528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3830_ack_0, ack => zeropad3D_F_CP_8333_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_3339/merge_stmt_3829_PhiAck/phi_stmt_3837_ack
      -- 
    phi_stmt_3837_ack_9529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3837_ack_0, ack => zeropad3D_F_CP_8333_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_3339/merge_stmt_3829_PhiAck/phi_stmt_3843_ack
      -- 
    phi_stmt_3843_ack_9530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3843_ack_0, ack => zeropad3D_F_CP_8333_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	1 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_3339/merge_stmt_3829_PhiAck/$exit
      -- 
    zeropad3D_F_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_F_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_F_CP_8333_elements(135) & zeropad3D_F_CP_8333_elements(136) & zeropad3D_F_CP_8333_elements(137);
      gj_zeropad3D_F_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_F_CP_8333_elements(138), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_3423_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3485_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3620_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3703_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3728_wire : std_logic_vector(31 downto 0);
    signal R_idxprom136_3714_resized : std_logic_vector(13 downto 0);
    signal R_idxprom136_3714_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom141_3739_resized : std_logic_vector(13 downto 0);
    signal R_idxprom141_3739_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3631_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3631_scaled : std_logic_vector(13 downto 0);
    signal add108_3671 : std_logic_vector(31 downto 0);
    signal add117_3676 : std_logic_vector(31 downto 0);
    signal add127_3691 : std_logic_vector(31 downto 0);
    signal add133_3696 : std_logic_vector(31 downto 0);
    signal add146_3759 : std_logic_vector(31 downto 0);
    signal add154_3779 : std_logic_vector(15 downto 0);
    signal add164_3436 : std_logic_vector(31 downto 0);
    signal add181_3457 : std_logic_vector(31 downto 0);
    signal add79_3467 : std_logic_vector(31 downto 0);
    signal add90_3608 : std_logic_vector(31 downto 0);
    signal add96_3613 : std_logic_vector(31 downto 0);
    signal add_3462 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3632_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3632_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3632_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3632_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3632_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3632_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3715_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3715_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3715_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3715_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3715_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3715_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3740_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3740_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3740_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3740_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3740_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3740_root_address : std_logic_vector(13 downto 0);
    signal arrayidx137_3717 : std_logic_vector(31 downto 0);
    signal arrayidx142_3742 : std_logic_vector(31 downto 0);
    signal arrayidx_3634 : std_logic_vector(31 downto 0);
    signal call1_3345 : std_logic_vector(7 downto 0);
    signal call2_3348 : std_logic_vector(7 downto 0);
    signal call3_3351 : std_logic_vector(7 downto 0);
    signal call4_3354 : std_logic_vector(7 downto 0);
    signal call5_3357 : std_logic_vector(7 downto 0);
    signal call6_3360 : std_logic_vector(7 downto 0);
    signal call_3342 : std_logic_vector(7 downto 0);
    signal cmp149_3766 : std_logic_vector(0 downto 0);
    signal cmp165_3797 : std_logic_vector(0 downto 0);
    signal cmp182_3822 : std_logic_vector(0 downto 0);
    signal cmp63_3534 : std_logic_vector(0 downto 0);
    signal cmp70_3558 : std_logic_vector(0 downto 0);
    signal cmp70x_xnot_3564 : std_logic_vector(0 downto 0);
    signal cmp80_3571 : std_logic_vector(0 downto 0);
    signal cmp_3521 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_3527 : std_logic_vector(0 downto 0);
    signal conv100_3646 : std_logic_vector(31 downto 0);
    signal conv10_3375 : std_logic_vector(15 downto 0);
    signal conv110_3487 : std_logic_vector(31 downto 0);
    signal conv145_3753 : std_logic_vector(31 downto 0);
    signal conv159_3792 : std_logic_vector(31 downto 0);
    signal conv173_3817 : std_logic_vector(31 downto 0);
    signal conv175_3440 : std_logic_vector(31 downto 0);
    signal conv36_3385 : std_logic_vector(31 downto 0);
    signal conv38_3389 : std_logic_vector(31 downto 0);
    signal conv42_3393 : std_logic_vector(31 downto 0);
    signal conv44_3397 : std_logic_vector(31 downto 0);
    signal conv51_3514 : std_logic_vector(31 downto 0);
    signal conv53_3406 : std_logic_vector(31 downto 0);
    signal conv67_3551 : std_logic_vector(31 downto 0);
    signal conv84_3588 : std_logic_vector(31 downto 0);
    signal conv86_3410 : std_logic_vector(31 downto 0);
    signal conv88_3593 : std_logic_vector(31 downto 0);
    signal conv92_3425 : std_logic_vector(31 downto 0);
    signal conv_3365 : std_logic_vector(15 downto 0);
    signal div11_3381 : std_logic_vector(15 downto 0);
    signal div177_3452 : std_logic_vector(31 downto 0);
    signal div_3371 : std_logic_vector(15 downto 0);
    signal idxprom136_3710 : std_logic_vector(63 downto 0);
    signal idxprom141_3735 : std_logic_vector(63 downto 0);
    signal idxprom_3627 : std_logic_vector(63 downto 0);
    signal inc170_3801 : std_logic_vector(15 downto 0);
    signal inc170x_xix_x2_3806 : std_logic_vector(15 downto 0);
    signal inc_3787 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_3837 : std_logic_vector(15 downto 0);
    signal ix_x2_3497 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_3843 : std_logic_vector(15 downto 0);
    signal jx_x1_3503 : std_logic_vector(15 downto 0);
    signal jx_x2_3812 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_3830 : std_logic_vector(15 downto 0);
    signal kx_x1_3490 : std_logic_vector(15 downto 0);
    signal mul107_3656 : std_logic_vector(31 downto 0);
    signal mul116_3666 : std_logic_vector(31 downto 0);
    signal mul126_3681 : std_logic_vector(31 downto 0);
    signal mul132_3686 : std_logic_vector(31 downto 0);
    signal mul176_3446 : std_logic_vector(31 downto 0);
    signal mul45_3402 : std_logic_vector(31 downto 0);
    signal mul89_3598 : std_logic_vector(31 downto 0);
    signal mul95_3603 : std_logic_vector(31 downto 0);
    signal mul_3473 : std_logic_vector(31 downto 0);
    signal orx_xcond196_3576 : std_logic_vector(0 downto 0);
    signal orx_xcond_3539 : std_logic_vector(0 downto 0);
    signal ptr_deref_3636_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3636_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3636_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3636_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3636_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3636_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3720_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3720_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3720_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3720_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3720_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3744_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3744_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3744_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3744_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3744_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3744_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext195_3416 : std_logic_vector(31 downto 0);
    signal sext_3478 : std_logic_vector(31 downto 0);
    signal shl_3431 : std_logic_vector(31 downto 0);
    signal shr135_3705 : std_logic_vector(31 downto 0);
    signal shr140_3730 : std_logic_vector(31 downto 0);
    signal shr_3622 : std_logic_vector(31 downto 0);
    signal sub115_3661 : std_logic_vector(31 downto 0);
    signal sub_3651 : std_logic_vector(31 downto 0);
    signal tmp138_3721 : std_logic_vector(63 downto 0);
    signal type_cast_3369_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3379_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3414_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3419_wire : std_logic_vector(31 downto 0);
    signal type_cast_3422_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3444_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3450_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3471_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3481_wire : std_logic_vector(31 downto 0);
    signal type_cast_3484_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3494_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3496_wire : std_logic_vector(15 downto 0);
    signal type_cast_3500_wire : std_logic_vector(15 downto 0);
    signal type_cast_3502_wire : std_logic_vector(15 downto 0);
    signal type_cast_3506_wire : std_logic_vector(15 downto 0);
    signal type_cast_3508_wire : std_logic_vector(15 downto 0);
    signal type_cast_3512_wire : std_logic_vector(31 downto 0);
    signal type_cast_3517_wire : std_logic_vector(31 downto 0);
    signal type_cast_3519_wire : std_logic_vector(31 downto 0);
    signal type_cast_3525_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3530_wire : std_logic_vector(31 downto 0);
    signal type_cast_3532_wire : std_logic_vector(31 downto 0);
    signal type_cast_3549_wire : std_logic_vector(31 downto 0);
    signal type_cast_3554_wire : std_logic_vector(31 downto 0);
    signal type_cast_3556_wire : std_logic_vector(31 downto 0);
    signal type_cast_3562_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3567_wire : std_logic_vector(31 downto 0);
    signal type_cast_3569_wire : std_logic_vector(31 downto 0);
    signal type_cast_3586_wire : std_logic_vector(31 downto 0);
    signal type_cast_3591_wire : std_logic_vector(31 downto 0);
    signal type_cast_3616_wire : std_logic_vector(31 downto 0);
    signal type_cast_3619_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3625_wire : std_logic_vector(63 downto 0);
    signal type_cast_3638_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3644_wire : std_logic_vector(31 downto 0);
    signal type_cast_3699_wire : std_logic_vector(31 downto 0);
    signal type_cast_3702_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3708_wire : std_logic_vector(63 downto 0);
    signal type_cast_3724_wire : std_logic_vector(31 downto 0);
    signal type_cast_3727_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3733_wire : std_logic_vector(63 downto 0);
    signal type_cast_3751_wire : std_logic_vector(31 downto 0);
    signal type_cast_3757_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3762_wire : std_logic_vector(31 downto 0);
    signal type_cast_3764_wire : std_logic_vector(31 downto 0);
    signal type_cast_3777_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3785_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3790_wire : std_logic_vector(31 downto 0);
    signal type_cast_3815_wire : std_logic_vector(31 downto 0);
    signal type_cast_3833_wire : std_logic_vector(15 downto 0);
    signal type_cast_3836_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3840_wire : std_logic_vector(15 downto 0);
    signal type_cast_3842_wire : std_logic_vector(15 downto 0);
    signal type_cast_3846_wire : std_logic_vector(15 downto 0);
    signal type_cast_3848_wire : std_logic_vector(15 downto 0);
    signal type_cast_3855_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_3632_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3632_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3632_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3632_resized_base_address <= "00000000000000";
    array_obj_ref_3715_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3715_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3715_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3715_resized_base_address <= "00000000000000";
    array_obj_ref_3740_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3740_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3740_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3740_resized_base_address <= "00000000000000";
    ptr_deref_3636_word_offset_0 <= "00000000000000";
    ptr_deref_3720_word_offset_0 <= "00000000000000";
    ptr_deref_3744_word_offset_0 <= "00000000000000";
    type_cast_3369_wire_constant <= "0000000000000001";
    type_cast_3379_wire_constant <= "0000000000000001";
    type_cast_3414_wire_constant <= "00000000000000000000000000010000";
    type_cast_3422_wire_constant <= "00000000000000000000000000010000";
    type_cast_3429_wire_constant <= "00000000000000000000000000000001";
    type_cast_3444_wire_constant <= "00000000000000000000000000000011";
    type_cast_3450_wire_constant <= "00000000000000000000000000000010";
    type_cast_3471_wire_constant <= "00000000000000000000000000010000";
    type_cast_3484_wire_constant <= "00000000000000000000000000010000";
    type_cast_3494_wire_constant <= "0000000000000000";
    type_cast_3525_wire_constant <= "1";
    type_cast_3562_wire_constant <= "1";
    type_cast_3619_wire_constant <= "00000000000000000000000000000010";
    type_cast_3638_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3702_wire_constant <= "00000000000000000000000000000010";
    type_cast_3727_wire_constant <= "00000000000000000000000000000010";
    type_cast_3757_wire_constant <= "00000000000000000000000000000100";
    type_cast_3777_wire_constant <= "0000000000000100";
    type_cast_3785_wire_constant <= "0000000000000001";
    type_cast_3836_wire_constant <= "0000000000000000";
    type_cast_3855_wire_constant <= "00000001";
    phi_stmt_3490: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3494_wire_constant & type_cast_3496_wire;
      req <= phi_stmt_3490_req_0 & phi_stmt_3490_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3490",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3490_ack_0,
          idata => idata,
          odata => kx_x1_3490,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3490
    phi_stmt_3497: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3500_wire & type_cast_3502_wire;
      req <= phi_stmt_3497_req_0 & phi_stmt_3497_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3497",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3497_ack_0,
          idata => idata,
          odata => ix_x2_3497,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3497
    phi_stmt_3503: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3506_wire & type_cast_3508_wire;
      req <= phi_stmt_3503_req_0 & phi_stmt_3503_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3503",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3503_ack_0,
          idata => idata,
          odata => jx_x1_3503,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3503
    phi_stmt_3830: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3833_wire & type_cast_3836_wire_constant;
      req <= phi_stmt_3830_req_0 & phi_stmt_3830_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3830",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3830_ack_0,
          idata => idata,
          odata => kx_x0x_xph_3830,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3830
    phi_stmt_3837: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3840_wire & type_cast_3842_wire;
      req <= phi_stmt_3837_req_0 & phi_stmt_3837_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3837",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3837_ack_0,
          idata => idata,
          odata => ix_x1x_xph_3837,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3837
    phi_stmt_3843: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3846_wire & type_cast_3848_wire;
      req <= phi_stmt_3843_req_0 & phi_stmt_3843_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3843",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3843_ack_0,
          idata => idata,
          odata => jx_x0x_xph_3843,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3843
    -- flow-through select operator MUX_3811_inst
    jx_x2_3812 <= div_3371 when (cmp165_3797(0) /=  '0') else inc_3787;
    addr_of_3633_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3633_final_reg_req_0;
      addr_of_3633_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3633_final_reg_req_1;
      addr_of_3633_final_reg_ack_1<= rack(0);
      addr_of_3633_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3633_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3632_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3634,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3716_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3716_final_reg_req_0;
      addr_of_3716_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3716_final_reg_req_1;
      addr_of_3716_final_reg_ack_1<= rack(0);
      addr_of_3716_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3716_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3715_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx137_3717,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3741_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3741_final_reg_req_0;
      addr_of_3741_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3741_final_reg_req_1;
      addr_of_3741_final_reg_ack_1<= rack(0);
      addr_of_3741_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3741_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3740_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx142_3742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3364_inst_req_0;
      type_cast_3364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3364_inst_req_1;
      type_cast_3364_inst_ack_1<= rack(0);
      type_cast_3364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_3345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_3365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3374_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3374_inst_req_0;
      type_cast_3374_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3374_inst_req_1;
      type_cast_3374_inst_ack_1<= rack(0);
      type_cast_3374_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3374_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_3342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_3375,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3384_inst_req_0;
      type_cast_3384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3384_inst_req_1;
      type_cast_3384_inst_ack_1<= rack(0);
      type_cast_3384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_3348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_3385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3388_inst_req_0;
      type_cast_3388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3388_inst_req_1;
      type_cast_3388_inst_ack_1<= rack(0);
      type_cast_3388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_3345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_3389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3392_inst_req_0;
      type_cast_3392_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3392_inst_req_1;
      type_cast_3392_inst_ack_1<= rack(0);
      type_cast_3392_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3392_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_3357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_3393,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3396_inst_req_0;
      type_cast_3396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3396_inst_req_1;
      type_cast_3396_inst_ack_1<= rack(0);
      type_cast_3396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_3354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_3397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3405_inst_req_0;
      type_cast_3405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3405_inst_req_1;
      type_cast_3405_inst_ack_1<= rack(0);
      type_cast_3405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_3360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_3406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3409_inst_req_0;
      type_cast_3409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3409_inst_req_1;
      type_cast_3409_inst_ack_1<= rack(0);
      type_cast_3409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_3357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_3410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3419_inst
    process(sext195_3416) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext195_3416(31 downto 0);
      type_cast_3419_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3424_inst
    process(ASHR_i32_i32_3423_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3423_wire(31 downto 0);
      conv92_3425 <= tmp_var; -- 
    end process;
    type_cast_3439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3439_inst_req_0;
      type_cast_3439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3439_inst_req_1;
      type_cast_3439_inst_ack_1<= rack(0);
      type_cast_3439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_3342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv175_3440,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3481_inst
    process(sext_3478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_3478(31 downto 0);
      type_cast_3481_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3486_inst
    process(ASHR_i32_i32_3485_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3485_wire(31 downto 0);
      conv110_3487 <= tmp_var; -- 
    end process;
    type_cast_3496_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3496_inst_req_0;
      type_cast_3496_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3496_inst_req_1;
      type_cast_3496_inst_ack_1<= rack(0);
      type_cast_3496_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3496_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_3830,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3496_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3500_inst_req_0;
      type_cast_3500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3500_inst_req_1;
      type_cast_3500_inst_ack_1<= rack(0);
      type_cast_3500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_3837,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3500_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3502_inst_req_0;
      type_cast_3502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3502_inst_req_1;
      type_cast_3502_inst_ack_1<= rack(0);
      type_cast_3502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div11_3381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3502_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3506_inst_req_0;
      type_cast_3506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3506_inst_req_1;
      type_cast_3506_inst_ack_1<= rack(0);
      type_cast_3506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_3371,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3506_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3508_inst_req_0;
      type_cast_3508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3508_inst_req_1;
      type_cast_3508_inst_ack_1<= rack(0);
      type_cast_3508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_3843,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3513_inst_req_0;
      type_cast_3513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3513_inst_req_1;
      type_cast_3513_inst_ack_1<= rack(0);
      type_cast_3513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3512_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_3514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3517_inst
    process(conv51_3514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv51_3514(31 downto 0);
      type_cast_3517_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3519_inst
    process(conv53_3406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_3406(31 downto 0);
      type_cast_3519_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3530_inst
    process(conv51_3514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv51_3514(31 downto 0);
      type_cast_3530_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3532_inst
    process(add_3462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_3462(31 downto 0);
      type_cast_3532_wire <= tmp_var; -- 
    end process;
    type_cast_3550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3550_inst_req_0;
      type_cast_3550_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3550_inst_req_1;
      type_cast_3550_inst_ack_1<= rack(0);
      type_cast_3550_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3550_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3549_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_3551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3554_inst
    process(conv67_3551) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv67_3551(31 downto 0);
      type_cast_3554_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3556_inst
    process(conv53_3406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_3406(31 downto 0);
      type_cast_3556_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3567_inst
    process(conv67_3551) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv67_3551(31 downto 0);
      type_cast_3567_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3569_inst
    process(add79_3467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add79_3467(31 downto 0);
      type_cast_3569_wire <= tmp_var; -- 
    end process;
    type_cast_3587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3587_inst_req_0;
      type_cast_3587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3587_inst_req_1;
      type_cast_3587_inst_ack_1<= rack(0);
      type_cast_3587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3586_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_3588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3592_inst_req_0;
      type_cast_3592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3592_inst_req_1;
      type_cast_3592_inst_ack_1<= rack(0);
      type_cast_3592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3591_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3616_inst
    process(add96_3613) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add96_3613(31 downto 0);
      type_cast_3616_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3621_inst
    process(ASHR_i32_i32_3620_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3620_wire(31 downto 0);
      shr_3622 <= tmp_var; -- 
    end process;
    type_cast_3626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3626_inst_req_0;
      type_cast_3626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3626_inst_req_1;
      type_cast_3626_inst_ack_1<= rack(0);
      type_cast_3626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3625_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3645_inst_req_0;
      type_cast_3645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3645_inst_req_1;
      type_cast_3645_inst_ack_1<= rack(0);
      type_cast_3645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3644_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_3646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3699_inst
    process(add117_3676) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add117_3676(31 downto 0);
      type_cast_3699_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3704_inst
    process(ASHR_i32_i32_3703_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3703_wire(31 downto 0);
      shr135_3705 <= tmp_var; -- 
    end process;
    type_cast_3709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3709_inst_req_0;
      type_cast_3709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3709_inst_req_1;
      type_cast_3709_inst_ack_1<= rack(0);
      type_cast_3709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3708_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom136_3710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3724_inst
    process(add133_3696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add133_3696(31 downto 0);
      type_cast_3724_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3729_inst
    process(ASHR_i32_i32_3728_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3728_wire(31 downto 0);
      shr140_3730 <= tmp_var; -- 
    end process;
    type_cast_3734_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3734_inst_req_0;
      type_cast_3734_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3734_inst_req_1;
      type_cast_3734_inst_ack_1<= rack(0);
      type_cast_3734_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3734_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3733_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom141_3735,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3752_inst_req_0;
      type_cast_3752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3752_inst_req_1;
      type_cast_3752_inst_ack_1<= rack(0);
      type_cast_3752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3751_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_3753,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3762_inst
    process(add146_3759) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add146_3759(31 downto 0);
      type_cast_3762_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3764_inst
    process(conv36_3385) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_3385(31 downto 0);
      type_cast_3764_wire <= tmp_var; -- 
    end process;
    type_cast_3791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3791_inst_req_0;
      type_cast_3791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3791_inst_req_1;
      type_cast_3791_inst_ack_1<= rack(0);
      type_cast_3791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3790_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_3792,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3800_inst_req_0;
      type_cast_3800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3800_inst_req_1;
      type_cast_3800_inst_ack_1<= rack(0);
      type_cast_3800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp165_3797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc170_3801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3816_inst_req_0;
      type_cast_3816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3816_inst_req_1;
      type_cast_3816_inst_ack_1<= rack(0);
      type_cast_3816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3815_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_3817,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3833_inst_req_0;
      type_cast_3833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3833_inst_req_1;
      type_cast_3833_inst_ack_1<= rack(0);
      type_cast_3833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add154_3779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3833_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3840_inst_req_0;
      type_cast_3840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3840_inst_req_1;
      type_cast_3840_inst_ack_1<= rack(0);
      type_cast_3840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_3497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3840_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3842_inst_req_0;
      type_cast_3842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3842_inst_req_1;
      type_cast_3842_inst_ack_1<= rack(0);
      type_cast_3842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc170x_xix_x2_3806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3842_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3846_inst_req_0;
      type_cast_3846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3846_inst_req_1;
      type_cast_3846_inst_ack_1<= rack(0);
      type_cast_3846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_3503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3846_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3848_inst_req_0;
      type_cast_3848_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3848_inst_req_1;
      type_cast_3848_inst_ack_1<= rack(0);
      type_cast_3848_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3848_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_3812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3848_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_3632_index_1_rename
    process(R_idxprom_3631_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3631_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3631_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3632_index_1_resize
    process(idxprom_3627) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3627;
      ov := iv(13 downto 0);
      R_idxprom_3631_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3632_root_address_inst
    process(array_obj_ref_3632_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3632_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3632_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3715_index_1_rename
    process(R_idxprom136_3714_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom136_3714_resized;
      ov(13 downto 0) := iv;
      R_idxprom136_3714_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3715_index_1_resize
    process(idxprom136_3710) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom136_3710;
      ov := iv(13 downto 0);
      R_idxprom136_3714_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3715_root_address_inst
    process(array_obj_ref_3715_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3715_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3715_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3740_index_1_rename
    process(R_idxprom141_3739_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom141_3739_resized;
      ov(13 downto 0) := iv;
      R_idxprom141_3739_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3740_index_1_resize
    process(idxprom141_3735) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom141_3735;
      ov := iv(13 downto 0);
      R_idxprom141_3739_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3740_root_address_inst
    process(array_obj_ref_3740_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3740_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3740_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_addr_0
    process(ptr_deref_3636_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3636_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3636_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_base_resize
    process(arrayidx_3634) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3634;
      ov := iv(13 downto 0);
      ptr_deref_3636_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_gather_scatter
    process(type_cast_3638_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3638_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3636_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_root_address_inst
    process(ptr_deref_3636_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3636_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3636_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3720_addr_0
    process(ptr_deref_3720_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3720_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3720_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3720_base_resize
    process(arrayidx137_3717) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx137_3717;
      ov := iv(13 downto 0);
      ptr_deref_3720_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3720_gather_scatter
    process(ptr_deref_3720_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3720_data_0;
      ov(63 downto 0) := iv;
      tmp138_3721 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3720_root_address_inst
    process(ptr_deref_3720_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3720_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3720_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3744_addr_0
    process(ptr_deref_3744_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3744_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3744_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3744_base_resize
    process(arrayidx142_3742) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx142_3742;
      ov := iv(13 downto 0);
      ptr_deref_3744_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3744_gather_scatter
    process(tmp138_3721) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp138_3721;
      ov(63 downto 0) := iv;
      ptr_deref_3744_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3744_root_address_inst
    process(ptr_deref_3744_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3744_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3744_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3540_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_3539;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3540_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3540_branch_req_0,
          ack0 => if_stmt_3540_branch_ack_0,
          ack1 => if_stmt_3540_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3577_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond196_3576;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3577_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3577_branch_req_0,
          ack0 => if_stmt_3577_branch_ack_0,
          ack1 => if_stmt_3577_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3767_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp149_3766;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3767_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3767_branch_req_0,
          ack0 => if_stmt_3767_branch_ack_0,
          ack1 => if_stmt_3767_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3823_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp182_3822;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3823_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3823_branch_req_0,
          ack0 => if_stmt_3823_branch_ack_0,
          ack1 => if_stmt_3823_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3778_inst
    process(kx_x1_3490) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_3490, type_cast_3777_wire_constant, tmp_var);
      add154_3779 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3786_inst
    process(jx_x1_3503) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_3503, type_cast_3785_wire_constant, tmp_var);
      inc_3787 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3805_inst
    process(inc170_3801, ix_x2_3497) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc170_3801, ix_x2_3497, tmp_var);
      inc170x_xix_x2_3806 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3435_inst
    process(shl_3431, conv38_3389) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_3431, conv38_3389, tmp_var);
      add164_3436 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3456_inst
    process(shl_3431, div177_3452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_3431, div177_3452, tmp_var);
      add181_3457 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3461_inst
    process(conv53_3406, div177_3452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv53_3406, div177_3452, tmp_var);
      add_3462 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3466_inst
    process(conv53_3406, conv38_3389) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv53_3406, conv38_3389, tmp_var);
      add79_3467 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3607_inst
    process(mul95_3603, conv84_3588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul95_3603, conv84_3588, tmp_var);
      add90_3608 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3612_inst
    process(add90_3608, mul89_3598) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add90_3608, mul89_3598, tmp_var);
      add96_3613 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3670_inst
    process(mul116_3666, conv100_3646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul116_3666, conv100_3646, tmp_var);
      add108_3671 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3675_inst
    process(add108_3671, mul107_3656) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add108_3671, mul107_3656, tmp_var);
      add117_3676 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3690_inst
    process(mul132_3686, conv100_3646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul132_3686, conv100_3646, tmp_var);
      add127_3691 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3695_inst
    process(add127_3691, mul126_3681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add127_3691, mul126_3681, tmp_var);
      add133_3696 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3758_inst
    process(conv145_3753) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv145_3753, type_cast_3757_wire_constant, tmp_var);
      add146_3759 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3538_inst
    process(cmpx_xnot_3527, cmp63_3534) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_3527, cmp63_3534, tmp_var);
      orx_xcond_3539 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3575_inst
    process(cmp70x_xnot_3564, cmp80_3571) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp70x_xnot_3564, cmp80_3571, tmp_var);
      orx_xcond196_3576 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3423_inst
    process(type_cast_3419_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3419_wire, type_cast_3422_wire_constant, tmp_var);
      ASHR_i32_i32_3423_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3485_inst
    process(type_cast_3481_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3481_wire, type_cast_3484_wire_constant, tmp_var);
      ASHR_i32_i32_3485_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3620_inst
    process(type_cast_3616_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3616_wire, type_cast_3619_wire_constant, tmp_var);
      ASHR_i32_i32_3620_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3703_inst
    process(type_cast_3699_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3699_wire, type_cast_3702_wire_constant, tmp_var);
      ASHR_i32_i32_3703_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3728_inst
    process(type_cast_3724_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3724_wire, type_cast_3727_wire_constant, tmp_var);
      ASHR_i32_i32_3728_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3796_inst
    process(conv159_3792, add164_3436) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv159_3792, add164_3436, tmp_var);
      cmp165_3797 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3821_inst
    process(conv173_3817, add181_3457) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv173_3817, add181_3457, tmp_var);
      cmp182_3822 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3370_inst
    process(conv_3365) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_3365, type_cast_3369_wire_constant, tmp_var);
      div_3371 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3380_inst
    process(conv10_3375) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv10_3375, type_cast_3379_wire_constant, tmp_var);
      div11_3381 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3451_inst
    process(mul176_3446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul176_3446, type_cast_3450_wire_constant, tmp_var);
      div177_3452 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3401_inst
    process(conv42_3393, conv44_3397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_3393, conv44_3397, tmp_var);
      mul45_3402 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3445_inst
    process(conv175_3440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv175_3440, type_cast_3444_wire_constant, tmp_var);
      mul176_3446 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3477_inst
    process(mul_3473, conv36_3385) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_3473, conv36_3385, tmp_var);
      sext_3478 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3597_inst
    process(conv88_3593, conv86_3410) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv88_3593, conv86_3410, tmp_var);
      mul89_3598 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3602_inst
    process(conv51_3514, conv92_3425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv51_3514, conv92_3425, tmp_var);
      mul95_3603 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3655_inst
    process(sub_3651, conv36_3385) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_3651, conv36_3385, tmp_var);
      mul107_3656 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3665_inst
    process(sub115_3661, conv110_3487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub115_3661, conv110_3487, tmp_var);
      mul116_3666 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3680_inst
    process(conv67_3551, conv86_3410) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv67_3551, conv86_3410, tmp_var);
      mul126_3681 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3685_inst
    process(conv51_3514, conv92_3425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv51_3514, conv92_3425, tmp_var);
      mul132_3686 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3415_inst
    process(mul45_3402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul45_3402, type_cast_3414_wire_constant, tmp_var);
      sext195_3416 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3430_inst
    process(conv53_3406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_3406, type_cast_3429_wire_constant, tmp_var);
      shl_3431 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3472_inst
    process(conv38_3389) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv38_3389, type_cast_3471_wire_constant, tmp_var);
      mul_3473 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3520_inst
    process(type_cast_3517_wire, type_cast_3519_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3517_wire, type_cast_3519_wire, tmp_var);
      cmp_3521 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3533_inst
    process(type_cast_3530_wire, type_cast_3532_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3530_wire, type_cast_3532_wire, tmp_var);
      cmp63_3534 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3557_inst
    process(type_cast_3554_wire, type_cast_3556_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3554_wire, type_cast_3556_wire, tmp_var);
      cmp70_3558 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3570_inst
    process(type_cast_3567_wire, type_cast_3569_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3567_wire, type_cast_3569_wire, tmp_var);
      cmp80_3571 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3765_inst
    process(type_cast_3762_wire, type_cast_3764_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3762_wire, type_cast_3764_wire, tmp_var);
      cmp149_3766 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3650_inst
    process(conv67_3551, conv53_3406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv67_3551, conv53_3406, tmp_var);
      sub_3651 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3660_inst
    process(conv51_3514, conv53_3406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv51_3514, conv53_3406, tmp_var);
      sub115_3661 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3526_inst
    process(cmp_3521) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_3521, type_cast_3525_wire_constant, tmp_var);
      cmpx_xnot_3527 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3563_inst
    process(cmp70_3558) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp70_3558, type_cast_3562_wire_constant, tmp_var);
      cmp70x_xnot_3564 <= tmp_var; --
    end process;
    -- shared split operator group (47) : array_obj_ref_3632_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3631_scaled;
      array_obj_ref_3632_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3632_index_offset_req_0;
      array_obj_ref_3632_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3632_index_offset_req_1;
      array_obj_ref_3632_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_3715_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom136_3714_scaled;
      array_obj_ref_3715_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3715_index_offset_req_0;
      array_obj_ref_3715_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3715_index_offset_req_1;
      array_obj_ref_3715_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : array_obj_ref_3740_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom141_3739_scaled;
      array_obj_ref_3740_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3740_index_offset_req_0;
      array_obj_ref_3740_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3740_index_offset_req_1;
      array_obj_ref_3740_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- unary operator type_cast_3512_inst
    process(ix_x2_3497) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_3497, tmp_var);
      type_cast_3512_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3549_inst
    process(jx_x1_3503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_3503, tmp_var);
      type_cast_3549_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3586_inst
    process(kx_x1_3490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_3490, tmp_var);
      type_cast_3586_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3591_inst
    process(jx_x1_3503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_3503, tmp_var);
      type_cast_3591_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3625_inst
    process(shr_3622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3622, tmp_var);
      type_cast_3625_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3644_inst
    process(kx_x1_3490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_3490, tmp_var);
      type_cast_3644_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3708_inst
    process(shr135_3705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr135_3705, tmp_var);
      type_cast_3708_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3733_inst
    process(shr140_3730) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr140_3730, tmp_var);
      type_cast_3733_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3751_inst
    process(kx_x1_3490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_3490, tmp_var);
      type_cast_3751_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3790_inst
    process(inc_3787) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3787, tmp_var);
      type_cast_3790_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3815_inst
    process(inc170x_xix_x2_3806) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc170x_xix_x2_3806, tmp_var);
      type_cast_3815_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_3720_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3720_load_0_req_0;
      ptr_deref_3720_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3720_load_0_req_1;
      ptr_deref_3720_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3720_word_address_0;
      ptr_deref_3720_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3636_store_0 ptr_deref_3744_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3636_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3744_store_0_req_0;
      ptr_deref_3636_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3744_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3636_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3744_store_0_req_1;
      ptr_deref_3636_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3744_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3636_word_address_0 & ptr_deref_3744_word_address_0;
      data_in <= ptr_deref_3636_data_0 & ptr_deref_3744_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block5_starting_3341_inst RPIPE_Block5_starting_3344_inst RPIPE_Block5_starting_3347_inst RPIPE_Block5_starting_3350_inst RPIPE_Block5_starting_3353_inst RPIPE_Block5_starting_3356_inst RPIPE_Block5_starting_3359_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block5_starting_3341_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block5_starting_3344_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block5_starting_3347_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block5_starting_3350_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block5_starting_3353_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block5_starting_3356_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block5_starting_3359_inst_req_0;
      RPIPE_Block5_starting_3341_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block5_starting_3344_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block5_starting_3347_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block5_starting_3350_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block5_starting_3353_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block5_starting_3356_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block5_starting_3359_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block5_starting_3341_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block5_starting_3344_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block5_starting_3347_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block5_starting_3350_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block5_starting_3353_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block5_starting_3356_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block5_starting_3359_inst_req_1;
      RPIPE_Block5_starting_3341_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block5_starting_3344_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block5_starting_3347_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block5_starting_3350_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block5_starting_3353_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block5_starting_3356_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block5_starting_3359_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call_3342 <= data_out(55 downto 48);
      call1_3345 <= data_out(47 downto 40);
      call2_3348 <= data_out(39 downto 32);
      call3_3351 <= data_out(31 downto 24);
      call4_3354 <= data_out(23 downto 16);
      call5_3357 <= data_out(15 downto 8);
      call6_3360 <= data_out(7 downto 0);
      Block5_starting_read_0_gI: SplitGuardInterface generic map(name => "Block5_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block5_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block5_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block5_starting_pipe_read_req(0),
          oack => Block5_starting_pipe_read_ack(0),
          odata => Block5_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block5_complete_3853_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block5_complete_3853_inst_req_0;
      WPIPE_Block5_complete_3853_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block5_complete_3853_inst_req_1;
      WPIPE_Block5_complete_3853_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_3855_wire_constant;
      Block5_complete_write_0_gI: SplitGuardInterface generic map(name => "Block5_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block5_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block5_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block5_complete_pipe_write_req(0),
          oack => Block5_complete_pipe_write_ack(0),
          odata => Block5_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_F_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_G is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block6_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block6_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block6_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block6_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block6_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block6_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_G;
architecture zeropad3D_G_arch of zeropad3D_G is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_G_CP_9547_start: Boolean;
  signal zeropad3D_G_CP_9547_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_3903_inst_ack_1 : boolean;
  signal type_cast_3903_inst_req_1 : boolean;
  signal type_cast_4064_inst_req_0 : boolean;
  signal type_cast_4027_inst_ack_0 : boolean;
  signal type_cast_4101_inst_ack_1 : boolean;
  signal type_cast_3907_inst_req_0 : boolean;
  signal type_cast_4106_inst_req_0 : boolean;
  signal type_cast_4140_inst_ack_1 : boolean;
  signal if_stmt_4054_branch_ack_1 : boolean;
  signal type_cast_3907_inst_ack_0 : boolean;
  signal type_cast_4106_inst_req_1 : boolean;
  signal type_cast_4106_inst_ack_1 : boolean;
  signal array_obj_ref_4146_index_offset_req_0 : boolean;
  signal array_obj_ref_4146_index_offset_ack_0 : boolean;
  signal array_obj_ref_4146_index_offset_req_1 : boolean;
  signal array_obj_ref_4146_index_offset_ack_1 : boolean;
  signal type_cast_4027_inst_req_0 : boolean;
  signal type_cast_3911_inst_ack_1 : boolean;
  signal type_cast_3964_inst_req_0 : boolean;
  signal if_stmt_4091_branch_req_0 : boolean;
  signal type_cast_3928_inst_ack_1 : boolean;
  signal type_cast_3964_inst_ack_0 : boolean;
  signal addr_of_4147_final_reg_req_0 : boolean;
  signal addr_of_4147_final_reg_ack_0 : boolean;
  signal addr_of_4147_final_reg_req_1 : boolean;
  signal addr_of_4147_final_reg_ack_1 : boolean;
  signal if_stmt_4054_branch_ack_0 : boolean;
  signal type_cast_3915_inst_req_1 : boolean;
  signal type_cast_4106_inst_ack_0 : boolean;
  signal type_cast_3915_inst_ack_1 : boolean;
  signal type_cast_3924_inst_req_1 : boolean;
  signal type_cast_3924_inst_ack_1 : boolean;
  signal type_cast_4101_inst_req_1 : boolean;
  signal if_stmt_4091_branch_ack_0 : boolean;
  signal type_cast_3911_inst_req_0 : boolean;
  signal type_cast_3911_inst_ack_0 : boolean;
  signal type_cast_3964_inst_req_1 : boolean;
  signal type_cast_4064_inst_req_1 : boolean;
  signal type_cast_3907_inst_req_1 : boolean;
  signal type_cast_4064_inst_ack_0 : boolean;
  signal type_cast_3924_inst_req_0 : boolean;
  signal type_cast_4027_inst_req_1 : boolean;
  signal type_cast_3964_inst_ack_1 : boolean;
  signal if_stmt_4091_branch_ack_1 : boolean;
  signal type_cast_4159_inst_req_1 : boolean;
  signal type_cast_4159_inst_ack_1 : boolean;
  signal type_cast_3928_inst_req_1 : boolean;
  signal if_stmt_4054_branch_req_0 : boolean;
  signal ptr_deref_4150_store_0_req_1 : boolean;
  signal ptr_deref_4150_store_0_ack_1 : boolean;
  signal type_cast_4027_inst_ack_1 : boolean;
  signal type_cast_4159_inst_req_0 : boolean;
  signal type_cast_4159_inst_ack_0 : boolean;
  signal type_cast_3928_inst_ack_0 : boolean;
  signal type_cast_4140_inst_req_1 : boolean;
  signal type_cast_4101_inst_ack_0 : boolean;
  signal type_cast_4140_inst_ack_0 : boolean;
  signal type_cast_4140_inst_req_0 : boolean;
  signal type_cast_4101_inst_req_0 : boolean;
  signal ptr_deref_4150_store_0_req_0 : boolean;
  signal ptr_deref_4150_store_0_ack_0 : boolean;
  signal type_cast_4064_inst_ack_1 : boolean;
  signal type_cast_3915_inst_ack_0 : boolean;
  signal type_cast_3924_inst_ack_0 : boolean;
  signal type_cast_3928_inst_req_0 : boolean;
  signal type_cast_3915_inst_req_0 : boolean;
  signal type_cast_3907_inst_ack_1 : boolean;
  signal type_cast_3911_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3864_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3864_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3864_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3864_inst_ack_1 : boolean;
  signal RPIPE_Block6_starting_3867_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3867_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3867_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3867_inst_ack_1 : boolean;
  signal RPIPE_Block6_starting_3870_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3870_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3870_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3870_inst_ack_1 : boolean;
  signal RPIPE_Block6_starting_3873_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3873_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3873_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3873_inst_ack_1 : boolean;
  signal RPIPE_Block6_starting_3876_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3876_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3876_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3876_inst_ack_1 : boolean;
  signal RPIPE_Block6_starting_3879_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3879_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3879_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3879_inst_ack_1 : boolean;
  signal RPIPE_Block6_starting_3882_inst_req_0 : boolean;
  signal RPIPE_Block6_starting_3882_inst_ack_0 : boolean;
  signal RPIPE_Block6_starting_3882_inst_req_1 : boolean;
  signal RPIPE_Block6_starting_3882_inst_ack_1 : boolean;
  signal type_cast_3887_inst_req_0 : boolean;
  signal type_cast_3887_inst_ack_0 : boolean;
  signal type_cast_3887_inst_req_1 : boolean;
  signal type_cast_3887_inst_ack_1 : boolean;
  signal type_cast_3903_inst_req_0 : boolean;
  signal type_cast_3903_inst_ack_0 : boolean;
  signal type_cast_4223_inst_req_0 : boolean;
  signal type_cast_4223_inst_ack_0 : boolean;
  signal type_cast_4223_inst_req_1 : boolean;
  signal type_cast_4223_inst_ack_1 : boolean;
  signal array_obj_ref_4229_index_offset_req_0 : boolean;
  signal array_obj_ref_4229_index_offset_ack_0 : boolean;
  signal array_obj_ref_4229_index_offset_req_1 : boolean;
  signal array_obj_ref_4229_index_offset_ack_1 : boolean;
  signal addr_of_4230_final_reg_req_0 : boolean;
  signal addr_of_4230_final_reg_ack_0 : boolean;
  signal addr_of_4230_final_reg_req_1 : boolean;
  signal addr_of_4230_final_reg_ack_1 : boolean;
  signal ptr_deref_4234_load_0_req_0 : boolean;
  signal ptr_deref_4234_load_0_ack_0 : boolean;
  signal ptr_deref_4234_load_0_req_1 : boolean;
  signal ptr_deref_4234_load_0_ack_1 : boolean;
  signal type_cast_4248_inst_req_0 : boolean;
  signal type_cast_4248_inst_ack_0 : boolean;
  signal type_cast_4248_inst_req_1 : boolean;
  signal type_cast_4248_inst_ack_1 : boolean;
  signal array_obj_ref_4254_index_offset_req_0 : boolean;
  signal array_obj_ref_4254_index_offset_ack_0 : boolean;
  signal array_obj_ref_4254_index_offset_req_1 : boolean;
  signal array_obj_ref_4254_index_offset_ack_1 : boolean;
  signal addr_of_4255_final_reg_req_0 : boolean;
  signal addr_of_4255_final_reg_ack_0 : boolean;
  signal addr_of_4255_final_reg_req_1 : boolean;
  signal addr_of_4255_final_reg_ack_1 : boolean;
  signal ptr_deref_4258_store_0_req_0 : boolean;
  signal ptr_deref_4258_store_0_ack_0 : boolean;
  signal ptr_deref_4258_store_0_req_1 : boolean;
  signal ptr_deref_4258_store_0_ack_1 : boolean;
  signal type_cast_4266_inst_req_0 : boolean;
  signal type_cast_4266_inst_ack_0 : boolean;
  signal type_cast_4266_inst_req_1 : boolean;
  signal type_cast_4266_inst_ack_1 : boolean;
  signal if_stmt_4281_branch_req_0 : boolean;
  signal if_stmt_4281_branch_ack_1 : boolean;
  signal if_stmt_4281_branch_ack_0 : boolean;
  signal type_cast_4305_inst_req_0 : boolean;
  signal type_cast_4305_inst_ack_0 : boolean;
  signal type_cast_4305_inst_req_1 : boolean;
  signal type_cast_4305_inst_ack_1 : boolean;
  signal type_cast_4314_inst_req_0 : boolean;
  signal type_cast_4314_inst_ack_0 : boolean;
  signal type_cast_4314_inst_req_1 : boolean;
  signal type_cast_4314_inst_ack_1 : boolean;
  signal type_cast_4331_inst_req_0 : boolean;
  signal type_cast_4331_inst_ack_0 : boolean;
  signal type_cast_4331_inst_req_1 : boolean;
  signal type_cast_4331_inst_ack_1 : boolean;
  signal if_stmt_4338_branch_req_0 : boolean;
  signal if_stmt_4338_branch_ack_1 : boolean;
  signal if_stmt_4338_branch_ack_0 : boolean;
  signal WPIPE_Block6_complete_4368_inst_req_0 : boolean;
  signal WPIPE_Block6_complete_4368_inst_ack_0 : boolean;
  signal WPIPE_Block6_complete_4368_inst_req_1 : boolean;
  signal WPIPE_Block6_complete_4368_inst_ack_1 : boolean;
  signal phi_stmt_4003_req_0 : boolean;
  signal type_cast_4013_inst_req_0 : boolean;
  signal type_cast_4013_inst_ack_0 : boolean;
  signal type_cast_4013_inst_req_1 : boolean;
  signal type_cast_4013_inst_ack_1 : boolean;
  signal phi_stmt_4010_req_0 : boolean;
  signal phi_stmt_4016_req_0 : boolean;
  signal type_cast_4009_inst_req_0 : boolean;
  signal type_cast_4009_inst_ack_0 : boolean;
  signal type_cast_4009_inst_req_1 : boolean;
  signal type_cast_4009_inst_ack_1 : boolean;
  signal phi_stmt_4003_req_1 : boolean;
  signal type_cast_4015_inst_req_0 : boolean;
  signal type_cast_4015_inst_ack_0 : boolean;
  signal type_cast_4015_inst_req_1 : boolean;
  signal type_cast_4015_inst_ack_1 : boolean;
  signal phi_stmt_4010_req_1 : boolean;
  signal type_cast_4022_inst_req_0 : boolean;
  signal type_cast_4022_inst_ack_0 : boolean;
  signal type_cast_4022_inst_req_1 : boolean;
  signal type_cast_4022_inst_ack_1 : boolean;
  signal phi_stmt_4016_req_1 : boolean;
  signal phi_stmt_4003_ack_0 : boolean;
  signal phi_stmt_4010_ack_0 : boolean;
  signal phi_stmt_4016_ack_0 : boolean;
  signal phi_stmt_4345_req_1 : boolean;
  signal type_cast_4357_inst_req_0 : boolean;
  signal type_cast_4357_inst_ack_0 : boolean;
  signal type_cast_4357_inst_req_1 : boolean;
  signal type_cast_4357_inst_ack_1 : boolean;
  signal phi_stmt_4352_req_1 : boolean;
  signal type_cast_4363_inst_req_0 : boolean;
  signal type_cast_4363_inst_ack_0 : boolean;
  signal type_cast_4363_inst_req_1 : boolean;
  signal type_cast_4363_inst_ack_1 : boolean;
  signal phi_stmt_4358_req_1 : boolean;
  signal type_cast_4348_inst_req_0 : boolean;
  signal type_cast_4348_inst_ack_0 : boolean;
  signal type_cast_4348_inst_req_1 : boolean;
  signal type_cast_4348_inst_ack_1 : boolean;
  signal phi_stmt_4345_req_0 : boolean;
  signal type_cast_4355_inst_req_0 : boolean;
  signal type_cast_4355_inst_ack_0 : boolean;
  signal type_cast_4355_inst_req_1 : boolean;
  signal type_cast_4355_inst_ack_1 : boolean;
  signal phi_stmt_4352_req_0 : boolean;
  signal type_cast_4361_inst_req_0 : boolean;
  signal type_cast_4361_inst_ack_0 : boolean;
  signal type_cast_4361_inst_req_1 : boolean;
  signal type_cast_4361_inst_ack_1 : boolean;
  signal phi_stmt_4358_req_0 : boolean;
  signal phi_stmt_4345_ack_0 : boolean;
  signal phi_stmt_4352_ack_0 : boolean;
  signal phi_stmt_4358_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_G_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_G_CP_9547_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_G_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_G_CP_9547_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_G_CP_9547_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_G_CP_9547_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_G_CP_9547: Block -- control-path 
    signal zeropad3D_G_CP_9547_elements: BooleanArray(134 downto 0);
    -- 
  begin -- 
    zeropad3D_G_CP_9547_elements(0) <= zeropad3D_G_CP_9547_start;
    zeropad3D_G_CP_9547_symbol <= zeropad3D_G_CP_9547_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3862/$entry
      -- CP-element group 0: 	 branch_block_stmt_3862/branch_block_stmt_3862__entry__
      -- CP-element group 0: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883__entry__
      -- CP-element group 0: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/$entry
      -- CP-element group 0: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Sample/rr
      -- 
    rr_9613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(0), ack => RPIPE_Block6_starting_3864_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	134 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	102 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_3862/merge_stmt_4344__exit__
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Update/cr
      -- 
    rr_10449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(1), ack => type_cast_4009_inst_req_0); -- 
    cr_10454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(1), ack => type_cast_4009_inst_req_1); -- 
    rr_10472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(1), ack => type_cast_4015_inst_req_0); -- 
    cr_10477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(1), ack => type_cast_4015_inst_req_1); -- 
    rr_10495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(1), ack => type_cast_4022_inst_req_0); -- 
    cr_10500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(1), ack => type_cast_4022_inst_req_1); -- 
    zeropad3D_G_CP_9547_elements(1) <= zeropad3D_G_CP_9547_elements(134);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Update/cr
      -- 
    ra_9614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3864_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(2)); -- 
    cr_9618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(2), ack => RPIPE_Block6_starting_3864_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3864_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Sample/rr
      -- 
    ca_9619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3864_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(3)); -- 
    rr_9627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(3), ack => RPIPE_Block6_starting_3867_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_update_start_
      -- CP-element group 4: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Update/cr
      -- 
    ra_9628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3867_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(4)); -- 
    cr_9632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(4), ack => RPIPE_Block6_starting_3867_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3867_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Sample/rr
      -- 
    ca_9633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3867_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(5)); -- 
    rr_9641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(5), ack => RPIPE_Block6_starting_3870_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Update/cr
      -- 
    ra_9642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3870_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(6)); -- 
    cr_9646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(6), ack => RPIPE_Block6_starting_3870_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3870_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Sample/rr
      -- 
    ca_9647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3870_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(7)); -- 
    rr_9655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(7), ack => RPIPE_Block6_starting_3873_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_update_start_
      -- CP-element group 8: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Update/cr
      -- 
    ra_9656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3873_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(8)); -- 
    cr_9660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(8), ack => RPIPE_Block6_starting_3873_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3873_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Sample/rr
      -- 
    ca_9661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3873_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(9)); -- 
    rr_9669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(9), ack => RPIPE_Block6_starting_3876_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_update_start_
      -- CP-element group 10: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Update/cr
      -- 
    ra_9670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3876_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(10)); -- 
    cr_9674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(10), ack => RPIPE_Block6_starting_3876_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3876_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Sample/rr
      -- 
    ca_9675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3876_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(11)); -- 
    rr_9683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(11), ack => RPIPE_Block6_starting_3879_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_update_start_
      -- CP-element group 12: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Update/cr
      -- 
    ra_9684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3879_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(12)); -- 
    cr_9688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(12), ack => RPIPE_Block6_starting_3879_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3879_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Sample/rr
      -- 
    ca_9689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3879_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(13)); -- 
    rr_9697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(13), ack => RPIPE_Block6_starting_3882_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_update_start_
      -- CP-element group 14: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Update/cr
      -- 
    ra_9698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3882_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(14)); -- 
    cr_9702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(14), ack => RPIPE_Block6_starting_3882_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15:  members (55) 
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883__exit__
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000__entry__
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/$exit
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3865_to_assign_stmt_3883/RPIPE_Block6_starting_3882_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_update_start_
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Sample/rr
      -- 
    ca_9703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block6_starting_3882_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(15)); -- 
    cr_9733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3903_inst_req_1); -- 
    rr_9742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3907_inst_req_0); -- 
    rr_9812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3964_inst_req_0); -- 
    cr_9775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3915_inst_req_1); -- 
    cr_9789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3924_inst_req_1); -- 
    rr_9756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3911_inst_req_0); -- 
    cr_9817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3964_inst_req_1); -- 
    cr_9747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3907_inst_req_1); -- 
    rr_9784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3924_inst_req_0); -- 
    cr_9803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3928_inst_req_1); -- 
    rr_9798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3928_inst_req_0); -- 
    rr_9770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3915_inst_req_0); -- 
    cr_9761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3911_inst_req_1); -- 
    rr_9714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3887_inst_req_0); -- 
    cr_9719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3887_inst_req_1); -- 
    rr_9728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(15), ack => type_cast_3903_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Sample/ra
      -- 
    ra_9715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3887_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3887_Update/ca
      -- 
    ca_9720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3887_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Sample/ra
      -- 
    ra_9729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3903_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3903_update_completed_
      -- 
    ca_9734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3903_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Sample/$exit
      -- 
    ra_9743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3907_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3907_Update/ca
      -- 
    ca_9748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3907_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Sample/ra
      -- 
    ra_9757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3911_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3911_Update/$exit
      -- 
    ca_9762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3911_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Sample/$exit
      -- 
    ra_9771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3915_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3915_update_completed_
      -- 
    ca_9776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3915_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Sample/ra
      -- 
    ra_9785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3924_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3924_update_completed_
      -- 
    ca_9790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3924_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Sample/ra
      -- 
    ra_9799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3928_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3928_Update/$exit
      -- 
    ca_9804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3928_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Sample/ra
      -- 
    ra_9813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3964_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/type_cast_3964_Update/ca
      -- 
    ca_9818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3964_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	21 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	25 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: 	90 
    -- CP-element group 32: 	91 
    -- CP-element group 32: 	93 
    -- CP-element group 32:  members (16) 
      -- CP-element group 32: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000__exit__
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody
      -- CP-element group 32: 	 branch_block_stmt_3862/assign_stmt_3888_to_assign_stmt_4000/$exit
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4003/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4016/$entry
      -- CP-element group 32: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/$entry
      -- 
    rr_10415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(32), ack => type_cast_4013_inst_req_0); -- 
    cr_10420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(32), ack => type_cast_4013_inst_req_1); -- 
    zeropad3D_G_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(31) & zeropad3D_G_CP_9547_elements(17) & zeropad3D_G_CP_9547_elements(19) & zeropad3D_G_CP_9547_elements(21) & zeropad3D_G_CP_9547_elements(23) & zeropad3D_G_CP_9547_elements(25) & zeropad3D_G_CP_9547_elements(27) & zeropad3D_G_CP_9547_elements(29);
      gj_zeropad3D_G_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	109 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_sample_completed_
      -- 
    ra_9830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4027_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	109 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (13) 
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054_else_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/$exit
      -- CP-element group 34: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054_eval_test/branch_req
      -- CP-element group 34: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_3862/R_orx_xcond_4055_place
      -- CP-element group 34: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053__exit__
      -- CP-element group 34: 	 branch_block_stmt_3862/if_stmt_4054__entry__
      -- 
    ca_9835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4027_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(34)); -- 
    branch_req_9843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(34), ack => if_stmt_4054_branch_req_0); -- 
    -- CP-element group 35:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (18) 
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_3862/if_stmt_4054_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/$entry
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_update_start_
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_3862/if_stmt_4054_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_3862/whilex_xbody_lorx_xlhsx_xfalse59
      -- CP-element group 35: 	 branch_block_stmt_3862/merge_stmt_4060__exit__
      -- CP-element group 35: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090__entry__
      -- CP-element group 35: 	 branch_block_stmt_3862/whilex_xbody_lorx_xlhsx_xfalse59_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_3862/whilex_xbody_lorx_xlhsx_xfalse59_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_3862/merge_stmt_4060_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_3862/merge_stmt_4060_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_3862/merge_stmt_4060_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_3862/merge_stmt_4060_PhiAck/dummy
      -- 
    if_choice_transition_9848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4054_branch_ack_1, ack => zeropad3D_G_CP_9547_elements(35)); -- 
    rr_9865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(35), ack => type_cast_4064_inst_req_0); -- 
    cr_9870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(35), ack => type_cast_4064_inst_req_1); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	110 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_3862/whilex_xbody_ifx_xthen
      -- CP-element group 36: 	 branch_block_stmt_3862/if_stmt_4054_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_3862/if_stmt_4054_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_3862/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_3862/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_9852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4054_branch_ack_0, ack => zeropad3D_G_CP_9547_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Sample/ra
      -- 
    ra_9866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4064_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (13) 
      -- CP-element group 38: 	 branch_block_stmt_3862/R_orx_xcond190_4092_place
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091_eval_test/branch_req
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091_if_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/$exit
      -- CP-element group 38: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091_else_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090/type_cast_4064_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_3862/assign_stmt_4065_to_assign_stmt_4090__exit__
      -- CP-element group 38: 	 branch_block_stmt_3862/if_stmt_4091__entry__
      -- 
    ca_9871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4064_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(38)); -- 
    branch_req_9879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(38), ack => if_stmt_4091_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_3862/lorx_xlhsx_xfalse59_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_3862/if_stmt_4091_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_3862/if_stmt_4091_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/merge_stmt_4155__exit__
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260__entry__
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_complete/req
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_complete/req
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_update_start_
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_3862/lorx_xlhsx_xfalse59_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/lorx_xlhsx_xfalse59_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_3862/merge_stmt_4155_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_3862/merge_stmt_4155_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_3862/merge_stmt_4155_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_3862/merge_stmt_4155_PhiAck/dummy
      -- 
    if_choice_transition_9884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4091_branch_ack_1, ack => zeropad3D_G_CP_9547_elements(39)); -- 
    cr_10047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => type_cast_4159_inst_req_1); -- 
    rr_10042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => type_cast_4159_inst_req_0); -- 
    cr_10061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => type_cast_4223_inst_req_1); -- 
    req_10092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => array_obj_ref_4229_index_offset_req_1); -- 
    req_10107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => addr_of_4230_final_reg_req_1); -- 
    cr_10152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => ptr_deref_4234_load_0_req_1); -- 
    cr_10171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => type_cast_4248_inst_req_1); -- 
    req_10202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => array_obj_ref_4254_index_offset_req_1); -- 
    req_10217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => addr_of_4255_final_reg_req_1); -- 
    cr_10267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(39), ack => ptr_deref_4258_store_0_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	110 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_3862/lorx_xlhsx_xfalse59_ifx_xthen
      -- CP-element group 40: 	 branch_block_stmt_3862/if_stmt_4091_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_3862/if_stmt_4091_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_3862/lorx_xlhsx_xfalse59_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_3862/lorx_xlhsx_xfalse59_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_9888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4091_branch_ack_0, ack => zeropad3D_G_CP_9547_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	110 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Sample/$exit
      -- 
    ra_9902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4101_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	110 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_update_completed_
      -- 
    ca_9907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4101_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	110 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Sample/ra
      -- 
    ra_9916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4106_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_update_completed_
      -- 
    ca_9921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4106_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Sample/$entry
      -- 
    rr_9929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(45), ack => type_cast_4140_inst_req_0); -- 
    zeropad3D_G_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(44) & zeropad3D_G_CP_9547_elements(42);
      gj_zeropad3D_G_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Sample/$exit
      -- 
    ra_9930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4140_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	110 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_computed_1
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Update/$exit
      -- 
    ca_9935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4140_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(47)); -- 
    req_9960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(47), ack => array_obj_ref_4146_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Sample/ack
      -- 
    ack_9961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4146_index_offset_ack_0, ack => zeropad3D_G_CP_9547_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	110 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_request/req
      -- CP-element group 49: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_root_address_calculated
      -- 
    ack_9966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4146_index_offset_ack_1, ack => zeropad3D_G_CP_9547_elements(49)); -- 
    req_9975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(49), ack => addr_of_4147_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_request/$exit
      -- CP-element group 50: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_request/ack
      -- 
    ack_9976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4147_final_reg_ack_0, ack => zeropad3D_G_CP_9547_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	110 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_word_addrgen/$entry
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/ptr_deref_4150_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/ptr_deref_4150_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/ptr_deref_4150_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/ptr_deref_4150_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/word_access_start/word_0/rr
      -- CP-element group 51: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/word_access_start/word_0/$entry
      -- 
    ack_9981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4147_final_reg_ack_1, ack => zeropad3D_G_CP_9547_elements(51)); -- 
    rr_10019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(51), ack => ptr_deref_4150_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/word_access_start/word_0/ra
      -- CP-element group 52: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Sample/word_access_start/word_0/$exit
      -- 
    ra_10020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4150_store_0_ack_0, ack => zeropad3D_G_CP_9547_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	110 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/word_access_complete/word_0/$exit
      -- 
    ca_10031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4150_store_0_ack_1, ack => zeropad3D_G_CP_9547_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: 	48 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	111 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/$exit
      -- CP-element group 54: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153__exit__
      -- CP-element group 54: 	 branch_block_stmt_3862/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_3862/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_3862/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_G_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(53) & zeropad3D_G_CP_9547_elements(48);
      gj_zeropad3D_G_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_sample_completed_
      -- 
    ra_10043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4159_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4159_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Sample/rr
      -- 
    ca_10048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4159_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(56)); -- 
    rr_10056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(56), ack => type_cast_4223_inst_req_0); -- 
    rr_10166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(56), ack => type_cast_4248_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Sample/ra
      -- 
    ra_10057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4223_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4223_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Sample/req
      -- 
    ca_10062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4223_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(58)); -- 
    req_10087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(58), ack => array_obj_ref_4229_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Sample/ack
      -- 
    ack_10088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4229_index_offset_ack_0, ack => zeropad3D_G_CP_9547_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4229_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_request/req
      -- 
    ack_10093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4229_index_offset_ack_1, ack => zeropad3D_G_CP_9547_elements(60)); -- 
    req_10102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(60), ack => addr_of_4230_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_request/ack
      -- 
    ack_10103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4230_final_reg_ack_0, ack => zeropad3D_G_CP_9547_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4230_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/word_access_start/word_0/rr
      -- 
    ack_10108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4230_final_reg_ack_1, ack => zeropad3D_G_CP_9547_elements(62)); -- 
    rr_10141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(62), ack => ptr_deref_4234_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Sample/word_access_start/word_0/ra
      -- 
    ra_10142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4234_load_0_ack_0, ack => zeropad3D_G_CP_9547_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/ptr_deref_4234_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/ptr_deref_4234_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/ptr_deref_4234_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4234_Update/ptr_deref_4234_Merge/merge_ack
      -- 
    ca_10153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4234_load_0_ack_1, ack => zeropad3D_G_CP_9547_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Sample/ra
      -- 
    ra_10167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4248_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/type_cast_4248_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_computed_1
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Sample/req
      -- 
    ca_10172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4248_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(66)); -- 
    req_10197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(66), ack => array_obj_ref_4254_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Sample/ack
      -- 
    ack_10198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4254_index_offset_ack_0, ack => zeropad3D_G_CP_9547_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/array_obj_ref_4254_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_request/req
      -- 
    ack_10203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4254_index_offset_ack_1, ack => zeropad3D_G_CP_9547_elements(68)); -- 
    req_10212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(68), ack => addr_of_4255_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_request/ack
      -- 
    ack_10213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4255_final_reg_ack_0, ack => zeropad3D_G_CP_9547_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/addr_of_4255_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_word_addrgen/root_register_ack
      -- 
    ack_10218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4255_final_reg_ack_1, ack => zeropad3D_G_CP_9547_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/ptr_deref_4258_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/ptr_deref_4258_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/ptr_deref_4258_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/ptr_deref_4258_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/word_access_start/word_0/rr
      -- 
    rr_10256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(71), ack => ptr_deref_4258_store_0_req_0); -- 
    zeropad3D_G_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(64) & zeropad3D_G_CP_9547_elements(70);
      gj_zeropad3D_G_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Sample/word_access_start/word_0/ra
      -- 
    ra_10257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4258_store_0_ack_0, ack => zeropad3D_G_CP_9547_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/ptr_deref_4258_Update/word_access_complete/word_0/ca
      -- 
    ca_10268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4258_store_0_ack_1, ack => zeropad3D_G_CP_9547_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	111 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260/$exit
      -- CP-element group 74: 	 branch_block_stmt_3862/assign_stmt_4160_to_assign_stmt_4260__exit__
      -- CP-element group 74: 	 branch_block_stmt_3862/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_3862/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_3862/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_G_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(59) & zeropad3D_G_CP_9547_elements(67) & zeropad3D_G_CP_9547_elements(73);
      gj_zeropad3D_G_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	111 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Sample/ra
      -- 
    ra_10280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4266_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	111 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280__exit__
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281__entry__
      -- CP-element group 76: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/$exit
      -- CP-element group 76: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_3862/R_cmp144_4282_place
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_3862/if_stmt_4281_else_link/$entry
      -- 
    ca_10285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4266_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(76)); -- 
    branch_req_10293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(76), ack => if_stmt_4281_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	127 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_3862/merge_stmt_4287__exit__
      -- CP-element group 77: 	 branch_block_stmt_3862/assign_stmt_4293__entry__
      -- CP-element group 77: 	 branch_block_stmt_3862/assign_stmt_4293__exit__
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184
      -- CP-element group 77: 	 branch_block_stmt_3862/if_stmt_4281_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_3862/if_stmt_4281_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xend_ifx_xthen146
      -- CP-element group 77: 	 branch_block_stmt_3862/assign_stmt_4293/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/assign_stmt_4293/$exit
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xend_ifx_xthen146_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xend_ifx_xthen146_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_3862/merge_stmt_4287_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_3862/merge_stmt_4287_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/merge_stmt_4287_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_3862/merge_stmt_4287_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Update/cr
      -- 
    if_choice_transition_10298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4281_branch_ack_1, ack => zeropad3D_G_CP_9547_elements(77)); -- 
    rr_10655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(77), ack => type_cast_4348_inst_req_0); -- 
    cr_10660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(77), ack => type_cast_4348_inst_req_1); -- 
    rr_10678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(77), ack => type_cast_4355_inst_req_0); -- 
    cr_10683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(77), ack => type_cast_4355_inst_req_1); -- 
    rr_10701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(77), ack => type_cast_4361_inst_req_0); -- 
    cr_10706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(77), ack => type_cast_4361_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (24) 
      -- CP-element group 78: 	 branch_block_stmt_3862/merge_stmt_4295__exit__
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337__entry__
      -- CP-element group 78: 	 branch_block_stmt_3862/if_stmt_4281_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_3862/if_stmt_4281_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_3862/ifx_xend_ifx_xelse151
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_update_start_
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_update_start_
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_update_start_
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_3862/ifx_xend_ifx_xelse151_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/ifx_xend_ifx_xelse151_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_3862/merge_stmt_4295_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_3862/merge_stmt_4295_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_3862/merge_stmt_4295_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_3862/merge_stmt_4295_PhiAck/dummy
      -- 
    else_choice_transition_10302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4281_branch_ack_0, ack => zeropad3D_G_CP_9547_elements(78)); -- 
    rr_10318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(78), ack => type_cast_4305_inst_req_0); -- 
    cr_10323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(78), ack => type_cast_4305_inst_req_1); -- 
    cr_10337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(78), ack => type_cast_4314_inst_req_1); -- 
    cr_10351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(78), ack => type_cast_4331_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Sample/ra
      -- 
    ra_10319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4305_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4305_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Sample/rr
      -- 
    ca_10324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4305_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(80)); -- 
    rr_10332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(80), ack => type_cast_4314_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Sample/ra
      -- 
    ra_10333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4314_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4314_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Sample/rr
      -- 
    ca_10338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4314_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(82)); -- 
    rr_10346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(82), ack => type_cast_4331_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Sample/ra
      -- 
    ra_10347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4331_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(83)); -- 
    -- CP-element group 84:  branch  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (13) 
      -- CP-element group 84: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337__exit__
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338__entry__
      -- CP-element group 84: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/$exit
      -- CP-element group 84: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_3862/assign_stmt_4301_to_assign_stmt_4337/type_cast_4331_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_3862/R_cmp176_4339_place
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_3862/if_stmt_4338_else_link/$entry
      -- 
    ca_10352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4331_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(84)); -- 
    branch_req_10360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(84), ack => if_stmt_4338_branch_req_0); -- 
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_3862/merge_stmt_4366__exit__
      -- CP-element group 85: 	 branch_block_stmt_3862/assign_stmt_4371__entry__
      -- CP-element group 85: 	 branch_block_stmt_3862/if_stmt_4338_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_3862/if_stmt_4338_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_3862/ifx_xelse151_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_3862/assign_stmt_4371/$entry
      -- CP-element group 85: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_3862/ifx_xelse151_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_3862/ifx_xelse151_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_3862/merge_stmt_4366_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_3862/merge_stmt_4366_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_3862/merge_stmt_4366_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_3862/merge_stmt_4366_PhiAck/dummy
      -- 
    if_choice_transition_10365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4338_branch_ack_1, ack => zeropad3D_G_CP_9547_elements(85)); -- 
    req_10382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(85), ack => WPIPE_Block6_complete_4368_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	114 
    -- CP-element group 86: 	116 
    -- CP-element group 86: 	117 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_3862/if_stmt_4338_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_3862/if_stmt_4338_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4345/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Update/cr
      -- 
    else_choice_transition_10369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4338_branch_ack_0, ack => zeropad3D_G_CP_9547_elements(86)); -- 
    rr_10606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(86), ack => type_cast_4357_inst_req_0); -- 
    cr_10611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(86), ack => type_cast_4357_inst_req_1); -- 
    rr_10629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(86), ack => type_cast_4363_inst_req_0); -- 
    cr_10634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(86), ack => type_cast_4363_inst_req_1); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_update_start_
      -- CP-element group 87: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Update/req
      -- 
    ack_10383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_complete_4368_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(87)); -- 
    req_10387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(87), ack => WPIPE_Block6_complete_4368_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_3862/$exit
      -- CP-element group 88: 	 branch_block_stmt_3862/branch_block_stmt_3862__exit__
      -- CP-element group 88: 	 branch_block_stmt_3862/assign_stmt_4371__exit__
      -- CP-element group 88: 	 branch_block_stmt_3862/return__
      -- CP-element group 88: 	 branch_block_stmt_3862/merge_stmt_4373__exit__
      -- CP-element group 88: 	 branch_block_stmt_3862/assign_stmt_4371/$exit
      -- CP-element group 88: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_3862/assign_stmt_4371/WPIPE_Block6_complete_4368_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_3862/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_3862/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_3862/merge_stmt_4373_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_3862/merge_stmt_4373_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_3862/merge_stmt_4373_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_3862/merge_stmt_4373_PhiAck/dummy
      -- 
    ack_10388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block6_complete_4368_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(88)); -- 
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	94 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4003/$exit
      -- CP-element group 89: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4007_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_req
      -- 
    phi_stmt_4003_req_10399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4003_req_10399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(89), ack => phi_stmt_4003_req_0); -- 
    -- Element group zeropad3D_G_CP_9547_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_G_CP_9547_elements(32), ack => zeropad3D_G_CP_9547_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	32 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Sample/ra
      -- 
    ra_10416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4013_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/Update/ca
      -- 
    ca_10421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4013_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/$exit
      -- CP-element group 92: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/$exit
      -- CP-element group 92: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4013/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_req
      -- 
    phi_stmt_4010_req_10422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4010_req_10422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(92), ack => phi_stmt_4010_req_0); -- 
    zeropad3D_G_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(90) & zeropad3D_G_CP_9547_elements(91);
      gj_zeropad3D_G_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	32 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4016/$exit
      -- CP-element group 93: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4020_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_req
      -- 
    phi_stmt_4016_req_10430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4016_req_10430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(93), ack => phi_stmt_4016_req_0); -- 
    -- Element group zeropad3D_G_CP_9547_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => zeropad3D_G_CP_9547_elements(32), ack => zeropad3D_G_CP_9547_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	105 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_3862/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_G_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(89) & zeropad3D_G_CP_9547_elements(92) & zeropad3D_G_CP_9547_elements(93);
      gj_zeropad3D_G_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Sample/ra
      -- 
    ra_10450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4009_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/Update/ca
      -- 
    ca_10455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4009_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/$exit
      -- CP-element group 97: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/$exit
      -- CP-element group 97: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_sources/type_cast_4009/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4003/phi_stmt_4003_req
      -- 
    phi_stmt_4003_req_10456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4003_req_10456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(97), ack => phi_stmt_4003_req_1); -- 
    zeropad3D_G_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_G_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(95) & zeropad3D_G_CP_9547_elements(96);
      gj_zeropad3D_G_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Sample/ra
      -- 
    ra_10473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4015_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/Update/ca
      -- 
    ca_10478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4015_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/$exit
      -- CP-element group 100: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/$exit
      -- CP-element group 100: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_sources/type_cast_4015/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4010/phi_stmt_4010_req
      -- 
    phi_stmt_4010_req_10479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4010_req_10479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(100), ack => phi_stmt_4010_req_1); -- 
    zeropad3D_G_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(98) & zeropad3D_G_CP_9547_elements(99);
      gj_zeropad3D_G_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Sample/ra
      -- 
    ra_10496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4022_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/Update/ca
      -- 
    ca_10501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4022_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/$exit
      -- CP-element group 103: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/$exit
      -- CP-element group 103: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_sources/type_cast_4022/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_4016/phi_stmt_4016_req
      -- 
    phi_stmt_4016_req_10502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4016_req_10502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(103), ack => phi_stmt_4016_req_1); -- 
    zeropad3D_G_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(101) & zeropad3D_G_CP_9547_elements(102);
      gj_zeropad3D_G_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_3862/ifx_xend184_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_G_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(97) & zeropad3D_G_CP_9547_elements(100) & zeropad3D_G_CP_9547_elements(103);
      gj_zeropad3D_G_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  merge  fork  transition  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	94 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_3862/merge_stmt_4002_PhiReqMerge
      -- CP-element group 105: 	 branch_block_stmt_3862/merge_stmt_4002_PhiAck/$entry
      -- 
    zeropad3D_G_CP_9547_elements(105) <= OrReduce(zeropad3D_G_CP_9547_elements(94) & zeropad3D_G_CP_9547_elements(104));
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_3862/merge_stmt_4002_PhiAck/phi_stmt_4003_ack
      -- 
    phi_stmt_4003_ack_10507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4003_ack_0, ack => zeropad3D_G_CP_9547_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_3862/merge_stmt_4002_PhiAck/phi_stmt_4010_ack
      -- 
    phi_stmt_4010_ack_10508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4010_ack_0, ack => zeropad3D_G_CP_9547_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_3862/merge_stmt_4002_PhiAck/phi_stmt_4016_ack
      -- 
    phi_stmt_4016_ack_10509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4016_ack_0, ack => zeropad3D_G_CP_9547_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	34 
    -- CP-element group 109: 	33 
    -- CP-element group 109:  members (10) 
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/type_cast_4027_update_start_
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053/$entry
      -- CP-element group 109: 	 branch_block_stmt_3862/merge_stmt_4002__exit__
      -- CP-element group 109: 	 branch_block_stmt_3862/assign_stmt_4028_to_assign_stmt_4053__entry__
      -- CP-element group 109: 	 branch_block_stmt_3862/merge_stmt_4002_PhiAck/$exit
      -- 
    rr_9829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(109), ack => type_cast_4027_inst_req_0); -- 
    cr_9834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(109), ack => type_cast_4027_inst_req_1); -- 
    zeropad3D_G_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(106) & zeropad3D_G_CP_9547_elements(107) & zeropad3D_G_CP_9547_elements(108);
      gj_zeropad3D_G_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  merge  fork  transition  place  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	40 
    -- CP-element group 110: 	36 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	51 
    -- CP-element group 110: 	53 
    -- CP-element group 110: 	43 
    -- CP-element group 110: 	41 
    -- CP-element group 110: 	47 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	44 
    -- CP-element group 110: 	42 
    -- CP-element group 110:  members (33) 
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_update_start
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/array_obj_ref_4146_final_index_sum_regn_Update/req
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_update_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_complete/req
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_update_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4106_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/addr_of_4147_update_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_update_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_update_start_
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/word_access_complete/word_0/cr
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/word_access_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4140_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/type_cast_4101_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153/ptr_deref_4150_Update/word_access_complete/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/merge_stmt_4097__exit__
      -- CP-element group 110: 	 branch_block_stmt_3862/assign_stmt_4102_to_assign_stmt_4153__entry__
      -- CP-element group 110: 	 branch_block_stmt_3862/merge_stmt_4097_PhiReqMerge
      -- CP-element group 110: 	 branch_block_stmt_3862/merge_stmt_4097_PhiAck/$entry
      -- CP-element group 110: 	 branch_block_stmt_3862/merge_stmt_4097_PhiAck/$exit
      -- CP-element group 110: 	 branch_block_stmt_3862/merge_stmt_4097_PhiAck/dummy
      -- 
    rr_9915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => type_cast_4106_inst_req_0); -- 
    cr_9920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => type_cast_4106_inst_req_1); -- 
    req_9965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => array_obj_ref_4146_index_offset_req_1); -- 
    req_9980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => addr_of_4147_final_reg_req_1); -- 
    cr_9906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => type_cast_4101_inst_req_1); -- 
    cr_10030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => ptr_deref_4150_store_0_req_1); -- 
    cr_9934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => type_cast_4140_inst_req_1); -- 
    rr_9901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(110), ack => type_cast_4101_inst_req_0); -- 
    zeropad3D_G_CP_9547_elements(110) <= OrReduce(zeropad3D_G_CP_9547_elements(40) & zeropad3D_G_CP_9547_elements(36));
    -- CP-element group 111:  merge  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	54 
    -- CP-element group 111: 	74 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	75 
    -- CP-element group 111: 	76 
    -- CP-element group 111:  members (13) 
      -- CP-element group 111: 	 branch_block_stmt_3862/merge_stmt_4262__exit__
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280__entry__
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/$entry
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_update_start_
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_3862/assign_stmt_4267_to_assign_stmt_4280/type_cast_4266_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_3862/merge_stmt_4262_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_3862/merge_stmt_4262_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_3862/merge_stmt_4262_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_3862/merge_stmt_4262_PhiAck/dummy
      -- 
    rr_10279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(111), ack => type_cast_4266_inst_req_0); -- 
    cr_10284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(111), ack => type_cast_4266_inst_req_1); -- 
    zeropad3D_G_CP_9547_elements(111) <= OrReduce(zeropad3D_G_CP_9547_elements(54) & zeropad3D_G_CP_9547_elements(74));
    -- CP-element group 112:  transition  output  delay-element  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	119 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4345/$exit
      -- CP-element group 112: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/$exit
      -- CP-element group 112: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4351_konst_delay_trans
      -- CP-element group 112: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_req
      -- 
    phi_stmt_4345_req_10590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4345_req_10590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(112), ack => phi_stmt_4345_req_1); -- 
    -- Element group zeropad3D_G_CP_9547_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => zeropad3D_G_CP_9547_elements(86), ack => zeropad3D_G_CP_9547_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Sample/ra
      -- 
    ra_10607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4357_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	86 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/Update/ca
      -- 
    ca_10612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4357_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	119 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/$exit
      -- CP-element group 115: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/$exit
      -- CP-element group 115: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4357/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_req
      -- 
    phi_stmt_4352_req_10613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4352_req_10613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(115), ack => phi_stmt_4352_req_1); -- 
    zeropad3D_G_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(113) & zeropad3D_G_CP_9547_elements(114);
      gj_zeropad3D_G_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Sample/ra
      -- 
    ra_10630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4363_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	86 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/Update/ca
      -- 
    ca_10635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4363_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/$exit
      -- CP-element group 118: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/$exit
      -- CP-element group 118: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4363/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_req
      -- 
    phi_stmt_4358_req_10636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4358_req_10636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(118), ack => phi_stmt_4358_req_1); -- 
    zeropad3D_G_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(116) & zeropad3D_G_CP_9547_elements(117);
      gj_zeropad3D_G_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	112 
    -- CP-element group 119: 	115 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	130 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_3862/ifx_xelse151_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_G_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(112) & zeropad3D_G_CP_9547_elements(115) & zeropad3D_G_CP_9547_elements(118);
      gj_zeropad3D_G_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Sample/ra
      -- 
    ra_10656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4348_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/Update/ca
      -- 
    ca_10661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4348_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	129 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/$exit
      -- CP-element group 122: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/$exit
      -- CP-element group 122: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_sources/type_cast_4348/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4345/phi_stmt_4345_req
      -- 
    phi_stmt_4345_req_10662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4345_req_10662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(122), ack => phi_stmt_4345_req_0); -- 
    zeropad3D_G_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(120) & zeropad3D_G_CP_9547_elements(121);
      gj_zeropad3D_G_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/ra
      -- 
    ra_10679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4355_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/ca
      -- 
    ca_10684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4355_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/$exit
      -- CP-element group 125: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/$exit
      -- CP-element group 125: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4352/phi_stmt_4352_req
      -- 
    phi_stmt_4352_req_10685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4352_req_10685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(125), ack => phi_stmt_4352_req_0); -- 
    zeropad3D_G_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(123) & zeropad3D_G_CP_9547_elements(124);
      gj_zeropad3D_G_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Sample/ra
      -- 
    ra_10702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4361_inst_ack_0, ack => zeropad3D_G_CP_9547_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	77 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/Update/ca
      -- 
    ca_10707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4361_inst_ack_1, ack => zeropad3D_G_CP_9547_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/$exit
      -- CP-element group 128: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/$exit
      -- CP-element group 128: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_sources/type_cast_4361/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_4358/phi_stmt_4358_req
      -- 
    phi_stmt_4358_req_10708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4358_req_10708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_G_CP_9547_elements(128), ack => phi_stmt_4358_req_0); -- 
    zeropad3D_G_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(126) & zeropad3D_G_CP_9547_elements(127);
      gj_zeropad3D_G_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_3862/ifx_xthen146_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_G_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(122) & zeropad3D_G_CP_9547_elements(125) & zeropad3D_G_CP_9547_elements(128);
      gj_zeropad3D_G_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_3862/merge_stmt_4344_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_3862/merge_stmt_4344_PhiAck/$entry
      -- 
    zeropad3D_G_CP_9547_elements(130) <= OrReduce(zeropad3D_G_CP_9547_elements(119) & zeropad3D_G_CP_9547_elements(129));
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_3862/merge_stmt_4344_PhiAck/phi_stmt_4345_ack
      -- 
    phi_stmt_4345_ack_10713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4345_ack_0, ack => zeropad3D_G_CP_9547_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_3862/merge_stmt_4344_PhiAck/phi_stmt_4352_ack
      -- 
    phi_stmt_4352_ack_10714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4352_ack_0, ack => zeropad3D_G_CP_9547_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_3862/merge_stmt_4344_PhiAck/phi_stmt_4358_ack
      -- 
    phi_stmt_4358_ack_10715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4358_ack_0, ack => zeropad3D_G_CP_9547_elements(133)); -- 
    -- CP-element group 134:  join  transition  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	1 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_3862/merge_stmt_4344_PhiAck/$exit
      -- 
    zeropad3D_G_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_G_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_G_CP_9547_elements(131) & zeropad3D_G_CP_9547_elements(132) & zeropad3D_G_CP_9547_elements(133);
      gj_zeropad3D_G_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_G_CP_9547_elements(134), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_3942_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3998_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4134_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4217_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4242_wire : std_logic_vector(31 downto 0);
    signal R_idxprom131_4228_resized : std_logic_vector(13 downto 0);
    signal R_idxprom131_4228_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom136_4253_resized : std_logic_vector(13 downto 0);
    signal R_idxprom136_4253_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_4145_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_4145_scaled : std_logic_vector(13 downto 0);
    signal add103_4185 : std_logic_vector(31 downto 0);
    signal add112_4190 : std_logic_vector(31 downto 0);
    signal add122_4205 : std_logic_vector(31 downto 0);
    signal add128_4210 : std_logic_vector(31 downto 0);
    signal add141_4273 : std_logic_vector(31 downto 0);
    signal add149_4293 : std_logic_vector(15 downto 0);
    signal add160_3961 : std_logic_vector(31 downto 0);
    signal add175_3970 : std_logic_vector(31 downto 0);
    signal add74_3980 : std_logic_vector(31 downto 0);
    signal add85_4122 : std_logic_vector(31 downto 0);
    signal add91_4127 : std_logic_vector(31 downto 0);
    signal add_3975 : std_logic_vector(31 downto 0);
    signal array_obj_ref_4146_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4146_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4146_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4146_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4146_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4146_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4229_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4229_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4229_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4229_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4229_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4229_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4254_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4254_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4254_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4254_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4254_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4254_root_address : std_logic_vector(13 downto 0);
    signal arrayidx132_4231 : std_logic_vector(31 downto 0);
    signal arrayidx137_4256 : std_logic_vector(31 downto 0);
    signal arrayidx_4148 : std_logic_vector(31 downto 0);
    signal call1_3868 : std_logic_vector(7 downto 0);
    signal call2_3871 : std_logic_vector(7 downto 0);
    signal call3_3874 : std_logic_vector(7 downto 0);
    signal call4_3877 : std_logic_vector(7 downto 0);
    signal call5_3880 : std_logic_vector(7 downto 0);
    signal call6_3883 : std_logic_vector(7 downto 0);
    signal call_3865 : std_logic_vector(7 downto 0);
    signal cmp144_4280 : std_logic_vector(0 downto 0);
    signal cmp161_4311 : std_logic_vector(0 downto 0);
    signal cmp176_4337 : std_logic_vector(0 downto 0);
    signal cmp57_4048 : std_logic_vector(0 downto 0);
    signal cmp64_4072 : std_logic_vector(0 downto 0);
    signal cmp64x_xnot_4078 : std_logic_vector(0 downto 0);
    signal cmp75_4085 : std_logic_vector(0 downto 0);
    signal cmp_4035 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_4041 : std_logic_vector(0 downto 0);
    signal conv105_4000 : std_logic_vector(31 downto 0);
    signal conv140_4267 : std_logic_vector(31 downto 0);
    signal conv154_4306 : std_logic_vector(31 downto 0);
    signal conv169_4332 : std_logic_vector(31 downto 0);
    signal conv171_3965 : std_logic_vector(31 downto 0);
    signal conv31_3904 : std_logic_vector(31 downto 0);
    signal conv33_3908 : std_logic_vector(31 downto 0);
    signal conv38_3912 : std_logic_vector(31 downto 0);
    signal conv40_3916 : std_logic_vector(31 downto 0);
    signal conv47_4028 : std_logic_vector(31 downto 0);
    signal conv49_3925 : std_logic_vector(31 downto 0);
    signal conv61_4065 : std_logic_vector(31 downto 0);
    signal conv79_4102 : std_logic_vector(31 downto 0);
    signal conv81_3929 : std_logic_vector(31 downto 0);
    signal conv83_4107 : std_logic_vector(31 downto 0);
    signal conv87_3944 : std_logic_vector(31 downto 0);
    signal conv95_4160 : std_logic_vector(31 downto 0);
    signal conv_3888 : std_logic_vector(15 downto 0);
    signal div157_3950 : std_logic_vector(31 downto 0);
    signal div_3894 : std_logic_vector(15 downto 0);
    signal idxprom131_4224 : std_logic_vector(63 downto 0);
    signal idxprom136_4249 : std_logic_vector(63 downto 0);
    signal idxprom_4141 : std_logic_vector(63 downto 0);
    signal inc166_4315 : std_logic_vector(15 downto 0);
    signal inc166x_xix_x2_4320 : std_logic_vector(15 downto 0);
    signal inc_4301 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_4352 : std_logic_vector(15 downto 0);
    signal ix_x2_4010 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_4358 : std_logic_vector(15 downto 0);
    signal jx_x1_4016 : std_logic_vector(15 downto 0);
    signal jx_x2_4327 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_4345 : std_logic_vector(15 downto 0);
    signal kx_x1_4003 : std_logic_vector(15 downto 0);
    signal mul102_4170 : std_logic_vector(31 downto 0);
    signal mul111_4180 : std_logic_vector(31 downto 0);
    signal mul121_4195 : std_logic_vector(31 downto 0);
    signal mul127_4200 : std_logic_vector(31 downto 0);
    signal mul34_3986 : std_logic_vector(31 downto 0);
    signal mul41_3921 : std_logic_vector(31 downto 0);
    signal mul84_4112 : std_logic_vector(31 downto 0);
    signal mul90_4117 : std_logic_vector(31 downto 0);
    signal mul_3900 : std_logic_vector(15 downto 0);
    signal orx_xcond190_4090 : std_logic_vector(0 downto 0);
    signal orx_xcond_4053 : std_logic_vector(0 downto 0);
    signal ptr_deref_4150_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4150_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4150_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4150_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4150_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4150_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4234_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4234_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4234_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4234_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4234_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4258_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4258_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4258_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4258_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4258_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4258_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext189_3935 : std_logic_vector(31 downto 0);
    signal sext_3991 : std_logic_vector(31 downto 0);
    signal shl_3956 : std_logic_vector(31 downto 0);
    signal shr130_4219 : std_logic_vector(31 downto 0);
    signal shr135_4244 : std_logic_vector(31 downto 0);
    signal shr_4136 : std_logic_vector(31 downto 0);
    signal sub110_4175 : std_logic_vector(31 downto 0);
    signal sub_4165 : std_logic_vector(31 downto 0);
    signal tmp133_4235 : std_logic_vector(63 downto 0);
    signal type_cast_3892_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3898_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3933_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3938_wire : std_logic_vector(31 downto 0);
    signal type_cast_3941_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3948_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3954_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3984_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3994_wire : std_logic_vector(31 downto 0);
    signal type_cast_3997_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4007_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4009_wire : std_logic_vector(15 downto 0);
    signal type_cast_4013_wire : std_logic_vector(15 downto 0);
    signal type_cast_4015_wire : std_logic_vector(15 downto 0);
    signal type_cast_4020_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4022_wire : std_logic_vector(15 downto 0);
    signal type_cast_4026_wire : std_logic_vector(31 downto 0);
    signal type_cast_4031_wire : std_logic_vector(31 downto 0);
    signal type_cast_4033_wire : std_logic_vector(31 downto 0);
    signal type_cast_4039_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_4044_wire : std_logic_vector(31 downto 0);
    signal type_cast_4046_wire : std_logic_vector(31 downto 0);
    signal type_cast_4063_wire : std_logic_vector(31 downto 0);
    signal type_cast_4068_wire : std_logic_vector(31 downto 0);
    signal type_cast_4070_wire : std_logic_vector(31 downto 0);
    signal type_cast_4076_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_4081_wire : std_logic_vector(31 downto 0);
    signal type_cast_4083_wire : std_logic_vector(31 downto 0);
    signal type_cast_4100_wire : std_logic_vector(31 downto 0);
    signal type_cast_4105_wire : std_logic_vector(31 downto 0);
    signal type_cast_4130_wire : std_logic_vector(31 downto 0);
    signal type_cast_4133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4139_wire : std_logic_vector(63 downto 0);
    signal type_cast_4152_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_4158_wire : std_logic_vector(31 downto 0);
    signal type_cast_4213_wire : std_logic_vector(31 downto 0);
    signal type_cast_4216_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4222_wire : std_logic_vector(63 downto 0);
    signal type_cast_4238_wire : std_logic_vector(31 downto 0);
    signal type_cast_4241_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4247_wire : std_logic_vector(63 downto 0);
    signal type_cast_4265_wire : std_logic_vector(31 downto 0);
    signal type_cast_4271_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4276_wire : std_logic_vector(31 downto 0);
    signal type_cast_4278_wire : std_logic_vector(31 downto 0);
    signal type_cast_4291_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4299_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4304_wire : std_logic_vector(31 downto 0);
    signal type_cast_4324_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4330_wire : std_logic_vector(31 downto 0);
    signal type_cast_4348_wire : std_logic_vector(15 downto 0);
    signal type_cast_4351_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4355_wire : std_logic_vector(15 downto 0);
    signal type_cast_4357_wire : std_logic_vector(15 downto 0);
    signal type_cast_4361_wire : std_logic_vector(15 downto 0);
    signal type_cast_4363_wire : std_logic_vector(15 downto 0);
    signal type_cast_4370_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_4146_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4146_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4146_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4146_resized_base_address <= "00000000000000";
    array_obj_ref_4229_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4229_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4229_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4229_resized_base_address <= "00000000000000";
    array_obj_ref_4254_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4254_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4254_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4254_resized_base_address <= "00000000000000";
    ptr_deref_4150_word_offset_0 <= "00000000000000";
    ptr_deref_4234_word_offset_0 <= "00000000000000";
    ptr_deref_4258_word_offset_0 <= "00000000000000";
    type_cast_3892_wire_constant <= "0000000000000010";
    type_cast_3898_wire_constant <= "0000000000000011";
    type_cast_3933_wire_constant <= "00000000000000000000000000010000";
    type_cast_3941_wire_constant <= "00000000000000000000000000010000";
    type_cast_3948_wire_constant <= "00000000000000000000000000000001";
    type_cast_3954_wire_constant <= "00000000000000000000000000000001";
    type_cast_3984_wire_constant <= "00000000000000000000000000010000";
    type_cast_3997_wire_constant <= "00000000000000000000000000010000";
    type_cast_4007_wire_constant <= "0000000000000000";
    type_cast_4020_wire_constant <= "0000000000000000";
    type_cast_4039_wire_constant <= "1";
    type_cast_4076_wire_constant <= "1";
    type_cast_4133_wire_constant <= "00000000000000000000000000000010";
    type_cast_4152_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4216_wire_constant <= "00000000000000000000000000000010";
    type_cast_4241_wire_constant <= "00000000000000000000000000000010";
    type_cast_4271_wire_constant <= "00000000000000000000000000000100";
    type_cast_4291_wire_constant <= "0000000000000100";
    type_cast_4299_wire_constant <= "0000000000000001";
    type_cast_4324_wire_constant <= "0000000000000000";
    type_cast_4351_wire_constant <= "0000000000000000";
    type_cast_4370_wire_constant <= "00000001";
    phi_stmt_4003: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4007_wire_constant & type_cast_4009_wire;
      req <= phi_stmt_4003_req_0 & phi_stmt_4003_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4003",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4003_ack_0,
          idata => idata,
          odata => kx_x1_4003,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4003
    phi_stmt_4010: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4013_wire & type_cast_4015_wire;
      req <= phi_stmt_4010_req_0 & phi_stmt_4010_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4010",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4010_ack_0,
          idata => idata,
          odata => ix_x2_4010,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4010
    phi_stmt_4016: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4020_wire_constant & type_cast_4022_wire;
      req <= phi_stmt_4016_req_0 & phi_stmt_4016_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4016",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4016_ack_0,
          idata => idata,
          odata => jx_x1_4016,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4016
    phi_stmt_4345: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4348_wire & type_cast_4351_wire_constant;
      req <= phi_stmt_4345_req_0 & phi_stmt_4345_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4345",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4345_ack_0,
          idata => idata,
          odata => kx_x0x_xph_4345,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4345
    phi_stmt_4352: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4355_wire & type_cast_4357_wire;
      req <= phi_stmt_4352_req_0 & phi_stmt_4352_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4352",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4352_ack_0,
          idata => idata,
          odata => ix_x1x_xph_4352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4352
    phi_stmt_4358: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4361_wire & type_cast_4363_wire;
      req <= phi_stmt_4358_req_0 & phi_stmt_4358_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4358",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4358_ack_0,
          idata => idata,
          odata => jx_x0x_xph_4358,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4358
    -- flow-through select operator MUX_4326_inst
    jx_x2_4327 <= type_cast_4324_wire_constant when (cmp161_4311(0) /=  '0') else inc_4301;
    addr_of_4147_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4147_final_reg_req_0;
      addr_of_4147_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4147_final_reg_req_1;
      addr_of_4147_final_reg_ack_1<= rack(0);
      addr_of_4147_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4147_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4146_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_4148,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4230_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4230_final_reg_req_0;
      addr_of_4230_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4230_final_reg_req_1;
      addr_of_4230_final_reg_ack_1<= rack(0);
      addr_of_4230_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4230_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4229_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx132_4231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4255_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4255_final_reg_req_0;
      addr_of_4255_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4255_final_reg_req_1;
      addr_of_4255_final_reg_ack_1<= rack(0);
      addr_of_4255_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4255_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4254_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx137_4256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3887_inst_req_0;
      type_cast_3887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3887_inst_req_1;
      type_cast_3887_inst_ack_1<= rack(0);
      type_cast_3887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_3865,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_3888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3903_inst_req_0;
      type_cast_3903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3903_inst_req_1;
      type_cast_3903_inst_ack_1<= rack(0);
      type_cast_3903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_3871,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_3904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3907_inst_req_0;
      type_cast_3907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3907_inst_req_1;
      type_cast_3907_inst_ack_1<= rack(0);
      type_cast_3907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_3868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_3908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3911_inst_req_0;
      type_cast_3911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3911_inst_req_1;
      type_cast_3911_inst_ack_1<= rack(0);
      type_cast_3911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_3880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_3912,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3915_inst_req_0;
      type_cast_3915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3915_inst_req_1;
      type_cast_3915_inst_ack_1<= rack(0);
      type_cast_3915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_3877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_3916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3924_inst_req_0;
      type_cast_3924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3924_inst_req_1;
      type_cast_3924_inst_ack_1<= rack(0);
      type_cast_3924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_3883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_3925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3928_inst_req_0;
      type_cast_3928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3928_inst_req_1;
      type_cast_3928_inst_ack_1<= rack(0);
      type_cast_3928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_3880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_3929,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3938_inst
    process(sext189_3935) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext189_3935(31 downto 0);
      type_cast_3938_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3943_inst
    process(ASHR_i32_i32_3942_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3942_wire(31 downto 0);
      conv87_3944 <= tmp_var; -- 
    end process;
    type_cast_3964_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3964_inst_req_0;
      type_cast_3964_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3964_inst_req_1;
      type_cast_3964_inst_ack_1<= rack(0);
      type_cast_3964_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3964_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_3865,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_3965,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3994_inst
    process(sext_3991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_3991(31 downto 0);
      type_cast_3994_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3999_inst
    process(ASHR_i32_i32_3998_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3998_wire(31 downto 0);
      conv105_4000 <= tmp_var; -- 
    end process;
    type_cast_4009_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4009_inst_req_0;
      type_cast_4009_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4009_inst_req_1;
      type_cast_4009_inst_ack_1<= rack(0);
      type_cast_4009_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4009_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_4345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4009_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4013_inst_req_0;
      type_cast_4013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4013_inst_req_1;
      type_cast_4013_inst_ack_1<= rack(0);
      type_cast_4013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul_3900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4013_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4015_inst_req_0;
      type_cast_4015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4015_inst_req_1;
      type_cast_4015_inst_ack_1<= rack(0);
      type_cast_4015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_4352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4015_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4022_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4022_inst_req_0;
      type_cast_4022_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4022_inst_req_1;
      type_cast_4022_inst_ack_1<= rack(0);
      type_cast_4022_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4022_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_4358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4022_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4027_inst_req_0;
      type_cast_4027_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4027_inst_req_1;
      type_cast_4027_inst_ack_1<= rack(0);
      type_cast_4027_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4027_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4026_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_4028,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4031_inst
    process(conv47_4028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_4028(31 downto 0);
      type_cast_4031_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4033_inst
    process(conv49_3925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_3925(31 downto 0);
      type_cast_4033_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4044_inst
    process(conv47_4028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_4028(31 downto 0);
      type_cast_4044_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4046_inst
    process(add_3975) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_3975(31 downto 0);
      type_cast_4046_wire <= tmp_var; -- 
    end process;
    type_cast_4064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4064_inst_req_0;
      type_cast_4064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4064_inst_req_1;
      type_cast_4064_inst_ack_1<= rack(0);
      type_cast_4064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4063_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_4065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4068_inst
    process(conv61_4065) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv61_4065(31 downto 0);
      type_cast_4068_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4070_inst
    process(conv49_3925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_3925(31 downto 0);
      type_cast_4070_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4081_inst
    process(conv61_4065) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv61_4065(31 downto 0);
      type_cast_4081_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4083_inst
    process(add74_3980) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add74_3980(31 downto 0);
      type_cast_4083_wire <= tmp_var; -- 
    end process;
    type_cast_4101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4101_inst_req_0;
      type_cast_4101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4101_inst_req_1;
      type_cast_4101_inst_ack_1<= rack(0);
      type_cast_4101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4100_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_4102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4106_inst_req_0;
      type_cast_4106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4106_inst_req_1;
      type_cast_4106_inst_ack_1<= rack(0);
      type_cast_4106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4105_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_4107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4130_inst
    process(add91_4127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add91_4127(31 downto 0);
      type_cast_4130_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4135_inst
    process(ASHR_i32_i32_4134_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4134_wire(31 downto 0);
      shr_4136 <= tmp_var; -- 
    end process;
    type_cast_4140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4140_inst_req_0;
      type_cast_4140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4140_inst_req_1;
      type_cast_4140_inst_ack_1<= rack(0);
      type_cast_4140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4139_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_4141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4159_inst_req_0;
      type_cast_4159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4159_inst_req_1;
      type_cast_4159_inst_ack_1<= rack(0);
      type_cast_4159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4158_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_4160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4213_inst
    process(add112_4190) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add112_4190(31 downto 0);
      type_cast_4213_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4218_inst
    process(ASHR_i32_i32_4217_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4217_wire(31 downto 0);
      shr130_4219 <= tmp_var; -- 
    end process;
    type_cast_4223_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4223_inst_req_0;
      type_cast_4223_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4223_inst_req_1;
      type_cast_4223_inst_ack_1<= rack(0);
      type_cast_4223_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4223_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4222_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom131_4224,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4238_inst
    process(add128_4210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add128_4210(31 downto 0);
      type_cast_4238_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4243_inst
    process(ASHR_i32_i32_4242_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4242_wire(31 downto 0);
      shr135_4244 <= tmp_var; -- 
    end process;
    type_cast_4248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4248_inst_req_0;
      type_cast_4248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4248_inst_req_1;
      type_cast_4248_inst_ack_1<= rack(0);
      type_cast_4248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4247_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom136_4249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4266_inst_req_0;
      type_cast_4266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4266_inst_req_1;
      type_cast_4266_inst_ack_1<= rack(0);
      type_cast_4266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4265_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_4267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4276_inst
    process(add141_4273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add141_4273(31 downto 0);
      type_cast_4276_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4278_inst
    process(conv31_3904) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv31_3904(31 downto 0);
      type_cast_4278_wire <= tmp_var; -- 
    end process;
    type_cast_4305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4305_inst_req_0;
      type_cast_4305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4305_inst_req_1;
      type_cast_4305_inst_ack_1<= rack(0);
      type_cast_4305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4304_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_4306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4314_inst_req_0;
      type_cast_4314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4314_inst_req_1;
      type_cast_4314_inst_ack_1<= rack(0);
      type_cast_4314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp161_4311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc166_4315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4331_inst_req_0;
      type_cast_4331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4331_inst_req_1;
      type_cast_4331_inst_ack_1<= rack(0);
      type_cast_4331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4330_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv169_4332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4348_inst_req_0;
      type_cast_4348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4348_inst_req_1;
      type_cast_4348_inst_ack_1<= rack(0);
      type_cast_4348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add149_4293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4348_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4355_inst_req_0;
      type_cast_4355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4355_inst_req_1;
      type_cast_4355_inst_ack_1<= rack(0);
      type_cast_4355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_4010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4355_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4357_inst_req_0;
      type_cast_4357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4357_inst_req_1;
      type_cast_4357_inst_ack_1<= rack(0);
      type_cast_4357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc166x_xix_x2_4320,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4357_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4361_inst_req_0;
      type_cast_4361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4361_inst_req_1;
      type_cast_4361_inst_ack_1<= rack(0);
      type_cast_4361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_4016,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4361_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4363_inst_req_0;
      type_cast_4363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4363_inst_req_1;
      type_cast_4363_inst_ack_1<= rack(0);
      type_cast_4363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_4327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4363_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_4146_index_1_rename
    process(R_idxprom_4145_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_4145_resized;
      ov(13 downto 0) := iv;
      R_idxprom_4145_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4146_index_1_resize
    process(idxprom_4141) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_4141;
      ov := iv(13 downto 0);
      R_idxprom_4145_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4146_root_address_inst
    process(array_obj_ref_4146_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4146_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4146_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4229_index_1_rename
    process(R_idxprom131_4228_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom131_4228_resized;
      ov(13 downto 0) := iv;
      R_idxprom131_4228_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4229_index_1_resize
    process(idxprom131_4224) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom131_4224;
      ov := iv(13 downto 0);
      R_idxprom131_4228_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4229_root_address_inst
    process(array_obj_ref_4229_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4229_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4229_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4254_index_1_rename
    process(R_idxprom136_4253_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom136_4253_resized;
      ov(13 downto 0) := iv;
      R_idxprom136_4253_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4254_index_1_resize
    process(idxprom136_4249) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom136_4249;
      ov := iv(13 downto 0);
      R_idxprom136_4253_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4254_root_address_inst
    process(array_obj_ref_4254_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4254_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4254_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4150_addr_0
    process(ptr_deref_4150_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4150_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4150_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4150_base_resize
    process(arrayidx_4148) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_4148;
      ov := iv(13 downto 0);
      ptr_deref_4150_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4150_gather_scatter
    process(type_cast_4152_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_4152_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_4150_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4150_root_address_inst
    process(ptr_deref_4150_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4150_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4150_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4234_addr_0
    process(ptr_deref_4234_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4234_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4234_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4234_base_resize
    process(arrayidx132_4231) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx132_4231;
      ov := iv(13 downto 0);
      ptr_deref_4234_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4234_gather_scatter
    process(ptr_deref_4234_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4234_data_0;
      ov(63 downto 0) := iv;
      tmp133_4235 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4234_root_address_inst
    process(ptr_deref_4234_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4234_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4234_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4258_addr_0
    process(ptr_deref_4258_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4258_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4258_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4258_base_resize
    process(arrayidx137_4256) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx137_4256;
      ov := iv(13 downto 0);
      ptr_deref_4258_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4258_gather_scatter
    process(tmp133_4235) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp133_4235;
      ov(63 downto 0) := iv;
      ptr_deref_4258_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4258_root_address_inst
    process(ptr_deref_4258_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4258_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4258_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_4054_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_4053;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4054_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4054_branch_req_0,
          ack0 => if_stmt_4054_branch_ack_0,
          ack1 => if_stmt_4054_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4091_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond190_4090;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4091_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4091_branch_req_0,
          ack0 => if_stmt_4091_branch_ack_0,
          ack1 => if_stmt_4091_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4281_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp144_4280;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4281_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4281_branch_req_0,
          ack0 => if_stmt_4281_branch_ack_0,
          ack1 => if_stmt_4281_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4338_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp176_4337;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4338_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4338_branch_req_0,
          ack0 => if_stmt_4338_branch_ack_0,
          ack1 => if_stmt_4338_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_4292_inst
    process(kx_x1_4003) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_4003, type_cast_4291_wire_constant, tmp_var);
      add149_4293 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4300_inst
    process(jx_x1_4016) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_4016, type_cast_4299_wire_constant, tmp_var);
      inc_4301 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4319_inst
    process(inc166_4315, ix_x2_4010) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc166_4315, ix_x2_4010, tmp_var);
      inc166x_xix_x2_4320 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3960_inst
    process(shl_3956, div157_3950) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_3956, div157_3950, tmp_var);
      add160_3961 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3969_inst
    process(shl_3956, conv171_3965) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_3956, conv171_3965, tmp_var);
      add175_3970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3974_inst
    process(conv49_3925, conv171_3965) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv49_3925, conv171_3965, tmp_var);
      add_3975 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3979_inst
    process(conv49_3925, div157_3950) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv49_3925, div157_3950, tmp_var);
      add74_3980 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4121_inst
    process(mul90_4117, conv79_4102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul90_4117, conv79_4102, tmp_var);
      add85_4122 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4126_inst
    process(add85_4122, mul84_4112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add85_4122, mul84_4112, tmp_var);
      add91_4127 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4184_inst
    process(mul111_4180, conv95_4160) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul111_4180, conv95_4160, tmp_var);
      add103_4185 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4189_inst
    process(add103_4185, mul102_4170) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add103_4185, mul102_4170, tmp_var);
      add112_4190 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4204_inst
    process(mul127_4200, conv95_4160) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul127_4200, conv95_4160, tmp_var);
      add122_4205 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4209_inst
    process(add122_4205, mul121_4195) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add122_4205, mul121_4195, tmp_var);
      add128_4210 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4272_inst
    process(conv140_4267) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv140_4267, type_cast_4271_wire_constant, tmp_var);
      add141_4273 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_4052_inst
    process(cmpx_xnot_4041, cmp57_4048) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_4041, cmp57_4048, tmp_var);
      orx_xcond_4053 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_4089_inst
    process(cmp64x_xnot_4078, cmp75_4085) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp64x_xnot_4078, cmp75_4085, tmp_var);
      orx_xcond190_4090 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3942_inst
    process(type_cast_3938_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3938_wire, type_cast_3941_wire_constant, tmp_var);
      ASHR_i32_i32_3942_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3998_inst
    process(type_cast_3994_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3994_wire, type_cast_3997_wire_constant, tmp_var);
      ASHR_i32_i32_3998_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4134_inst
    process(type_cast_4130_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4130_wire, type_cast_4133_wire_constant, tmp_var);
      ASHR_i32_i32_4134_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4217_inst
    process(type_cast_4213_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4213_wire, type_cast_4216_wire_constant, tmp_var);
      ASHR_i32_i32_4217_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4242_inst
    process(type_cast_4238_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4238_wire, type_cast_4241_wire_constant, tmp_var);
      ASHR_i32_i32_4242_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4310_inst
    process(conv154_4306, add160_3961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv154_4306, add160_3961, tmp_var);
      cmp161_4311 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4336_inst
    process(conv169_4332, add175_3970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv169_4332, add175_3970, tmp_var);
      cmp176_4337 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3893_inst
    process(conv_3888) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_3888, type_cast_3892_wire_constant, tmp_var);
      div_3894 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3949_inst
    process(conv33_3908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv33_3908, type_cast_3948_wire_constant, tmp_var);
      div157_3950 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3899_inst
    process(div_3894) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(div_3894, type_cast_3898_wire_constant, tmp_var);
      mul_3900 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3920_inst
    process(conv38_3912, conv40_3916) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv38_3912, conv40_3916, tmp_var);
      mul41_3921 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3990_inst
    process(mul34_3986, conv31_3904) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul34_3986, conv31_3904, tmp_var);
      sext_3991 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4111_inst
    process(conv83_4107, conv81_3929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv83_4107, conv81_3929, tmp_var);
      mul84_4112 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4116_inst
    process(conv47_4028, conv87_3944) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv47_4028, conv87_3944, tmp_var);
      mul90_4117 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4169_inst
    process(sub_4165, conv31_3904) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_4165, conv31_3904, tmp_var);
      mul102_4170 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4179_inst
    process(sub110_4175, conv105_4000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub110_4175, conv105_4000, tmp_var);
      mul111_4180 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4194_inst
    process(conv61_4065, conv81_3929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv61_4065, conv81_3929, tmp_var);
      mul121_4195 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4199_inst
    process(conv47_4028, conv87_3944) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv47_4028, conv87_3944, tmp_var);
      mul127_4200 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3934_inst
    process(mul41_3921) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul41_3921, type_cast_3933_wire_constant, tmp_var);
      sext189_3935 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3955_inst
    process(conv49_3925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_3925, type_cast_3954_wire_constant, tmp_var);
      shl_3956 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3985_inst
    process(conv33_3908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv33_3908, type_cast_3984_wire_constant, tmp_var);
      mul34_3986 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4034_inst
    process(type_cast_4031_wire, type_cast_4033_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4031_wire, type_cast_4033_wire, tmp_var);
      cmp_4035 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4047_inst
    process(type_cast_4044_wire, type_cast_4046_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4044_wire, type_cast_4046_wire, tmp_var);
      cmp57_4048 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4071_inst
    process(type_cast_4068_wire, type_cast_4070_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4068_wire, type_cast_4070_wire, tmp_var);
      cmp64_4072 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4084_inst
    process(type_cast_4081_wire, type_cast_4083_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4081_wire, type_cast_4083_wire, tmp_var);
      cmp75_4085 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4279_inst
    process(type_cast_4276_wire, type_cast_4278_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4276_wire, type_cast_4278_wire, tmp_var);
      cmp144_4280 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4164_inst
    process(conv61_4065, conv49_3925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv61_4065, conv49_3925, tmp_var);
      sub_4165 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4174_inst
    process(conv47_4028, conv49_3925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv47_4028, conv49_3925, tmp_var);
      sub110_4175 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_4040_inst
    process(cmp_4035) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_4035, type_cast_4039_wire_constant, tmp_var);
      cmpx_xnot_4041 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_4077_inst
    process(cmp64_4072) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp64_4072, type_cast_4076_wire_constant, tmp_var);
      cmp64x_xnot_4078 <= tmp_var; --
    end process;
    -- shared split operator group (46) : array_obj_ref_4146_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_4145_scaled;
      array_obj_ref_4146_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4146_index_offset_req_0;
      array_obj_ref_4146_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4146_index_offset_req_1;
      array_obj_ref_4146_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_4229_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom131_4228_scaled;
      array_obj_ref_4229_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4229_index_offset_req_0;
      array_obj_ref_4229_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4229_index_offset_req_1;
      array_obj_ref_4229_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_4254_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom136_4253_scaled;
      array_obj_ref_4254_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4254_index_offset_req_0;
      array_obj_ref_4254_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4254_index_offset_req_1;
      array_obj_ref_4254_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- unary operator type_cast_4026_inst
    process(ix_x2_4010) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_4010, tmp_var);
      type_cast_4026_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4063_inst
    process(jx_x1_4016) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_4016, tmp_var);
      type_cast_4063_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4100_inst
    process(kx_x1_4003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_4003, tmp_var);
      type_cast_4100_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4105_inst
    process(jx_x1_4016) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_4016, tmp_var);
      type_cast_4105_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4139_inst
    process(shr_4136) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_4136, tmp_var);
      type_cast_4139_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4158_inst
    process(kx_x1_4003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_4003, tmp_var);
      type_cast_4158_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4222_inst
    process(shr130_4219) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr130_4219, tmp_var);
      type_cast_4222_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4247_inst
    process(shr135_4244) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr135_4244, tmp_var);
      type_cast_4247_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4265_inst
    process(kx_x1_4003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_4003, tmp_var);
      type_cast_4265_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4304_inst
    process(inc_4301) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_4301, tmp_var);
      type_cast_4304_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4330_inst
    process(inc166x_xix_x2_4320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc166x_xix_x2_4320, tmp_var);
      type_cast_4330_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_4234_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_4234_load_0_req_0;
      ptr_deref_4234_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_4234_load_0_req_1;
      ptr_deref_4234_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_4234_word_address_0;
      ptr_deref_4234_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_4258_store_0 ptr_deref_4150_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_4258_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4150_store_0_req_0;
      ptr_deref_4258_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4150_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_4258_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4150_store_0_req_1;
      ptr_deref_4258_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4150_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_4258_word_address_0 & ptr_deref_4150_word_address_0;
      data_in <= ptr_deref_4258_data_0 & ptr_deref_4150_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block6_starting_3882_inst RPIPE_Block6_starting_3879_inst RPIPE_Block6_starting_3876_inst RPIPE_Block6_starting_3873_inst RPIPE_Block6_starting_3870_inst RPIPE_Block6_starting_3867_inst RPIPE_Block6_starting_3864_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block6_starting_3882_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block6_starting_3879_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block6_starting_3876_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block6_starting_3873_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block6_starting_3870_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block6_starting_3867_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block6_starting_3864_inst_req_0;
      RPIPE_Block6_starting_3882_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block6_starting_3879_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block6_starting_3876_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block6_starting_3873_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block6_starting_3870_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block6_starting_3867_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block6_starting_3864_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block6_starting_3882_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block6_starting_3879_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block6_starting_3876_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block6_starting_3873_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block6_starting_3870_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block6_starting_3867_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block6_starting_3864_inst_req_1;
      RPIPE_Block6_starting_3882_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block6_starting_3879_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block6_starting_3876_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block6_starting_3873_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block6_starting_3870_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block6_starting_3867_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block6_starting_3864_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call6_3883 <= data_out(55 downto 48);
      call5_3880 <= data_out(47 downto 40);
      call4_3877 <= data_out(39 downto 32);
      call3_3874 <= data_out(31 downto 24);
      call2_3871 <= data_out(23 downto 16);
      call1_3868 <= data_out(15 downto 8);
      call_3865 <= data_out(7 downto 0);
      Block6_starting_read_0_gI: SplitGuardInterface generic map(name => "Block6_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block6_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block6_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block6_starting_pipe_read_req(0),
          oack => Block6_starting_pipe_read_ack(0),
          odata => Block6_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block6_complete_4368_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block6_complete_4368_inst_req_0;
      WPIPE_Block6_complete_4368_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block6_complete_4368_inst_req_1;
      WPIPE_Block6_complete_4368_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_4370_wire_constant;
      Block6_complete_write_0_gI: SplitGuardInterface generic map(name => "Block6_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block6_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block6_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block6_complete_pipe_write_req(0),
          oack => Block6_complete_pipe_write_ack(0),
          odata => Block6_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_G_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_H is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block7_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block7_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block7_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block7_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block7_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block7_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_H;
architecture zeropad3D_H_arch of zeropad3D_H is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_H_CP_10732_start: Boolean;
  signal zeropad3D_H_CP_10732_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block7_starting_4382_inst_req_1 : boolean;
  signal type_cast_4540_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4379_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4391_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4379_inst_ack_1 : boolean;
  signal RPIPE_Block7_starting_4382_inst_ack_1 : boolean;
  signal type_cast_4528_inst_ack_1 : boolean;
  signal RPIPE_Block7_starting_4382_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4385_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4385_inst_req_0 : boolean;
  signal RPIPE_Block7_starting_4388_inst_req_1 : boolean;
  signal type_cast_4534_inst_ack_1 : boolean;
  signal phi_stmt_4529_req_1 : boolean;
  signal RPIPE_Block7_starting_4379_inst_req_0 : boolean;
  signal RPIPE_Block7_starting_4388_inst_req_0 : boolean;
  signal RPIPE_Block7_starting_4388_inst_ack_0 : boolean;
  signal phi_stmt_4522_req_1 : boolean;
  signal type_cast_4540_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4385_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4391_inst_ack_1 : boolean;
  signal RPIPE_Block7_starting_4382_inst_req_0 : boolean;
  signal type_cast_4534_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4385_inst_ack_1 : boolean;
  signal RPIPE_Block7_starting_4379_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4394_inst_req_0 : boolean;
  signal RPIPE_Block7_starting_4394_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4391_inst_req_0 : boolean;
  signal RPIPE_Block7_starting_4391_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4394_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4388_inst_ack_1 : boolean;
  signal type_cast_4528_inst_req_1 : boolean;
  signal type_cast_4540_inst_req_0 : boolean;
  signal type_cast_4540_inst_ack_1 : boolean;
  signal phi_stmt_4875_ack_0 : boolean;
  signal type_cast_4868_inst_req_1 : boolean;
  signal type_cast_4868_inst_ack_1 : boolean;
  signal phi_stmt_4535_req_1 : boolean;
  signal phi_stmt_4862_ack_0 : boolean;
  signal phi_stmt_4869_ack_0 : boolean;
  signal phi_stmt_4869_req_0 : boolean;
  signal type_cast_4878_inst_req_0 : boolean;
  signal type_cast_4878_inst_ack_0 : boolean;
  signal type_cast_4874_inst_req_0 : boolean;
  signal type_cast_4868_inst_req_0 : boolean;
  signal type_cast_4868_inst_ack_0 : boolean;
  signal type_cast_4874_inst_ack_0 : boolean;
  signal type_cast_4872_inst_req_0 : boolean;
  signal phi_stmt_4522_ack_0 : boolean;
  signal type_cast_4872_inst_ack_0 : boolean;
  signal type_cast_4880_inst_req_0 : boolean;
  signal type_cast_4878_inst_req_1 : boolean;
  signal type_cast_4874_inst_req_1 : boolean;
  signal type_cast_4880_inst_ack_0 : boolean;
  signal type_cast_4878_inst_ack_1 : boolean;
  signal type_cast_4874_inst_ack_1 : boolean;
  signal phi_stmt_4875_req_0 : boolean;
  signal phi_stmt_4869_req_1 : boolean;
  signal phi_stmt_4862_req_1 : boolean;
  signal type_cast_4872_inst_req_1 : boolean;
  signal type_cast_4872_inst_ack_1 : boolean;
  signal RPIPE_Block7_starting_4394_inst_ack_1 : boolean;
  signal RPIPE_Block7_starting_4397_inst_req_0 : boolean;
  signal RPIPE_Block7_starting_4397_inst_ack_0 : boolean;
  signal RPIPE_Block7_starting_4397_inst_req_1 : boolean;
  signal RPIPE_Block7_starting_4397_inst_ack_1 : boolean;
  signal type_cast_4402_inst_req_0 : boolean;
  signal type_cast_4402_inst_ack_0 : boolean;
  signal type_cast_4402_inst_req_1 : boolean;
  signal type_cast_4402_inst_ack_1 : boolean;
  signal type_cast_4412_inst_req_0 : boolean;
  signal type_cast_4412_inst_ack_0 : boolean;
  signal type_cast_4412_inst_req_1 : boolean;
  signal type_cast_4412_inst_ack_1 : boolean;
  signal type_cast_4428_inst_req_0 : boolean;
  signal type_cast_4428_inst_ack_0 : boolean;
  signal type_cast_4428_inst_req_1 : boolean;
  signal type_cast_4428_inst_ack_1 : boolean;
  signal type_cast_4432_inst_req_0 : boolean;
  signal type_cast_4432_inst_ack_0 : boolean;
  signal type_cast_4432_inst_req_1 : boolean;
  signal type_cast_4432_inst_ack_1 : boolean;
  signal type_cast_4436_inst_req_0 : boolean;
  signal type_cast_4436_inst_ack_0 : boolean;
  signal type_cast_4436_inst_req_1 : boolean;
  signal type_cast_4436_inst_ack_1 : boolean;
  signal type_cast_4440_inst_req_0 : boolean;
  signal type_cast_4440_inst_ack_0 : boolean;
  signal type_cast_4440_inst_req_1 : boolean;
  signal type_cast_4440_inst_ack_1 : boolean;
  signal type_cast_4449_inst_req_0 : boolean;
  signal type_cast_4449_inst_ack_0 : boolean;
  signal type_cast_4449_inst_req_1 : boolean;
  signal type_cast_4449_inst_ack_1 : boolean;
  signal type_cast_4453_inst_req_0 : boolean;
  signal type_cast_4453_inst_ack_0 : boolean;
  signal type_cast_4453_inst_req_1 : boolean;
  signal type_cast_4453_inst_ack_1 : boolean;
  signal type_cast_4483_inst_req_0 : boolean;
  signal type_cast_4483_inst_ack_0 : boolean;
  signal type_cast_4483_inst_req_1 : boolean;
  signal type_cast_4483_inst_ack_1 : boolean;
  signal type_cast_4545_inst_req_0 : boolean;
  signal type_cast_4545_inst_ack_0 : boolean;
  signal type_cast_4545_inst_req_1 : boolean;
  signal type_cast_4545_inst_ack_1 : boolean;
  signal if_stmt_4572_branch_req_0 : boolean;
  signal if_stmt_4572_branch_ack_1 : boolean;
  signal if_stmt_4572_branch_ack_0 : boolean;
  signal type_cast_4582_inst_req_0 : boolean;
  signal type_cast_4582_inst_ack_0 : boolean;
  signal type_cast_4582_inst_req_1 : boolean;
  signal type_cast_4582_inst_ack_1 : boolean;
  signal if_stmt_4609_branch_req_0 : boolean;
  signal if_stmt_4609_branch_ack_1 : boolean;
  signal if_stmt_4609_branch_ack_0 : boolean;
  signal type_cast_4619_inst_req_0 : boolean;
  signal type_cast_4619_inst_ack_0 : boolean;
  signal type_cast_4619_inst_req_1 : boolean;
  signal type_cast_4619_inst_ack_1 : boolean;
  signal type_cast_4624_inst_req_0 : boolean;
  signal type_cast_4624_inst_ack_0 : boolean;
  signal type_cast_4624_inst_req_1 : boolean;
  signal type_cast_4624_inst_ack_1 : boolean;
  signal type_cast_4658_inst_req_0 : boolean;
  signal type_cast_4658_inst_ack_0 : boolean;
  signal type_cast_4658_inst_req_1 : boolean;
  signal type_cast_4658_inst_ack_1 : boolean;
  signal array_obj_ref_4664_index_offset_req_0 : boolean;
  signal array_obj_ref_4664_index_offset_ack_0 : boolean;
  signal array_obj_ref_4664_index_offset_req_1 : boolean;
  signal array_obj_ref_4664_index_offset_ack_1 : boolean;
  signal addr_of_4665_final_reg_req_0 : boolean;
  signal addr_of_4665_final_reg_ack_0 : boolean;
  signal addr_of_4665_final_reg_req_1 : boolean;
  signal addr_of_4665_final_reg_ack_1 : boolean;
  signal type_cast_4534_inst_ack_0 : boolean;
  signal type_cast_4534_inst_req_0 : boolean;
  signal phi_stmt_4535_ack_0 : boolean;
  signal ptr_deref_4668_store_0_req_0 : boolean;
  signal ptr_deref_4668_store_0_ack_0 : boolean;
  signal phi_stmt_4529_ack_0 : boolean;
  signal ptr_deref_4668_store_0_req_1 : boolean;
  signal ptr_deref_4668_store_0_ack_1 : boolean;
  signal phi_stmt_4862_req_0 : boolean;
  signal type_cast_4677_inst_req_0 : boolean;
  signal type_cast_4677_inst_ack_0 : boolean;
  signal type_cast_4677_inst_req_1 : boolean;
  signal type_cast_4677_inst_ack_1 : boolean;
  signal phi_stmt_4875_req_1 : boolean;
  signal type_cast_4741_inst_req_0 : boolean;
  signal type_cast_4741_inst_ack_0 : boolean;
  signal type_cast_4528_inst_ack_0 : boolean;
  signal type_cast_4741_inst_req_1 : boolean;
  signal type_cast_4741_inst_ack_1 : boolean;
  signal type_cast_4880_inst_ack_1 : boolean;
  signal type_cast_4880_inst_req_1 : boolean;
  signal array_obj_ref_4747_index_offset_req_0 : boolean;
  signal array_obj_ref_4747_index_offset_ack_0 : boolean;
  signal array_obj_ref_4747_index_offset_req_1 : boolean;
  signal array_obj_ref_4747_index_offset_ack_1 : boolean;
  signal addr_of_4748_final_reg_req_0 : boolean;
  signal addr_of_4748_final_reg_ack_0 : boolean;
  signal addr_of_4748_final_reg_req_1 : boolean;
  signal addr_of_4748_final_reg_ack_1 : boolean;
  signal ptr_deref_4752_load_0_req_0 : boolean;
  signal ptr_deref_4752_load_0_ack_0 : boolean;
  signal ptr_deref_4752_load_0_req_1 : boolean;
  signal ptr_deref_4752_load_0_ack_1 : boolean;
  signal type_cast_4766_inst_req_0 : boolean;
  signal type_cast_4766_inst_ack_0 : boolean;
  signal type_cast_4766_inst_req_1 : boolean;
  signal type_cast_4766_inst_ack_1 : boolean;
  signal array_obj_ref_4772_index_offset_req_0 : boolean;
  signal array_obj_ref_4772_index_offset_ack_0 : boolean;
  signal array_obj_ref_4772_index_offset_req_1 : boolean;
  signal array_obj_ref_4772_index_offset_ack_1 : boolean;
  signal addr_of_4773_final_reg_req_0 : boolean;
  signal addr_of_4773_final_reg_ack_0 : boolean;
  signal addr_of_4773_final_reg_req_1 : boolean;
  signal addr_of_4773_final_reg_ack_1 : boolean;
  signal ptr_deref_4776_store_0_req_0 : boolean;
  signal ptr_deref_4776_store_0_ack_0 : boolean;
  signal ptr_deref_4776_store_0_req_1 : boolean;
  signal ptr_deref_4776_store_0_ack_1 : boolean;
  signal type_cast_4784_inst_req_0 : boolean;
  signal type_cast_4784_inst_ack_0 : boolean;
  signal type_cast_4784_inst_req_1 : boolean;
  signal type_cast_4784_inst_ack_1 : boolean;
  signal if_stmt_4799_branch_req_0 : boolean;
  signal if_stmt_4799_branch_ack_1 : boolean;
  signal if_stmt_4799_branch_ack_0 : boolean;
  signal type_cast_4823_inst_req_0 : boolean;
  signal type_cast_4823_inst_ack_0 : boolean;
  signal type_cast_4823_inst_req_1 : boolean;
  signal type_cast_4823_inst_ack_1 : boolean;
  signal type_cast_4832_inst_req_0 : boolean;
  signal type_cast_4832_inst_ack_0 : boolean;
  signal type_cast_4832_inst_req_1 : boolean;
  signal type_cast_4832_inst_ack_1 : boolean;
  signal type_cast_4848_inst_req_0 : boolean;
  signal type_cast_4848_inst_ack_0 : boolean;
  signal type_cast_4848_inst_req_1 : boolean;
  signal type_cast_4848_inst_ack_1 : boolean;
  signal if_stmt_4855_branch_req_0 : boolean;
  signal if_stmt_4855_branch_ack_1 : boolean;
  signal if_stmt_4855_branch_ack_0 : boolean;
  signal WPIPE_Block7_complete_4885_inst_req_0 : boolean;
  signal WPIPE_Block7_complete_4885_inst_ack_0 : boolean;
  signal WPIPE_Block7_complete_4885_inst_req_1 : boolean;
  signal WPIPE_Block7_complete_4885_inst_ack_1 : boolean;
  signal phi_stmt_4522_req_0 : boolean;
  signal type_cast_4532_inst_req_0 : boolean;
  signal type_cast_4532_inst_ack_0 : boolean;
  signal type_cast_4532_inst_req_1 : boolean;
  signal type_cast_4532_inst_ack_1 : boolean;
  signal phi_stmt_4529_req_0 : boolean;
  signal type_cast_4538_inst_req_0 : boolean;
  signal type_cast_4538_inst_ack_0 : boolean;
  signal type_cast_4538_inst_req_1 : boolean;
  signal type_cast_4538_inst_ack_1 : boolean;
  signal phi_stmt_4535_req_0 : boolean;
  signal type_cast_4528_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_H_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_H_CP_10732_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_H_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_H_CP_10732_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_H_CP_10732_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_H_CP_10732_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_H_CP_10732: Block -- control-path 
    signal zeropad3D_H_CP_10732_elements: BooleanArray(138 downto 0);
    -- 
  begin -- 
    zeropad3D_H_CP_10732_elements(0) <= zeropad3D_H_CP_10732_start;
    zeropad3D_H_CP_10732_symbol <= zeropad3D_H_CP_10732_elements(90);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_4377/$entry
      -- CP-element group 0: 	 branch_block_stmt_4377/branch_block_stmt_4377__entry__
      -- CP-element group 0: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398__entry__
      -- 
    rr_10798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(0), ack => RPIPE_Block7_starting_4379_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	138 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	100 
    -- CP-element group 1: 	102 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	105 
    -- CP-element group 1: 	106 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/merge_stmt_4861__exit__
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Sample/rr
      -- 
    cr_11714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(1), ack => type_cast_4540_inst_req_1); -- 
    cr_11691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(1), ack => type_cast_4534_inst_req_1); -- 
    cr_11668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(1), ack => type_cast_4528_inst_req_1); -- 
    rr_11709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(1), ack => type_cast_4540_inst_req_0); -- 
    rr_11686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(1), ack => type_cast_4534_inst_req_0); -- 
    rr_11663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(1), ack => type_cast_4528_inst_req_0); -- 
    zeropad3D_H_CP_10732_elements(1) <= zeropad3D_H_CP_10732_elements(138);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_update_start_
      -- CP-element group 2: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Sample/ra
      -- 
    ra_10799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4379_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(2)); -- 
    cr_10803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(2), ack => RPIPE_Block7_starting_4379_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4379_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Sample/rr
      -- 
    ca_10804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4379_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(3)); -- 
    rr_10812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(3), ack => RPIPE_Block7_starting_4382_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_update_start_
      -- CP-element group 4: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_sample_completed_
      -- 
    ra_10813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4382_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(4)); -- 
    cr_10817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(4), ack => RPIPE_Block7_starting_4382_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4382_update_completed_
      -- 
    ca_10818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4382_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(5)); -- 
    rr_10826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(5), ack => RPIPE_Block7_starting_4385_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_update_start_
      -- CP-element group 6: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Sample/ra
      -- 
    ra_10827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4385_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(6)); -- 
    cr_10831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(6), ack => RPIPE_Block7_starting_4385_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4385_Update/ca
      -- 
    ca_10832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4385_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(7)); -- 
    rr_10840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(7), ack => RPIPE_Block7_starting_4388_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_update_start_
      -- CP-element group 8: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_sample_completed_
      -- 
    ra_10841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4388_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(8)); -- 
    cr_10845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(8), ack => RPIPE_Block7_starting_4388_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4388_Update/ca
      -- 
    ca_10846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4388_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(9)); -- 
    rr_10854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(9), ack => RPIPE_Block7_starting_4391_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_update_start_
      -- CP-element group 10: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Sample/ra
      -- 
    ra_10855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4391_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(10)); -- 
    cr_10859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(10), ack => RPIPE_Block7_starting_4391_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4391_Update/$exit
      -- 
    ca_10860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4391_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(11)); -- 
    rr_10868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(11), ack => RPIPE_Block7_starting_4394_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_update_start_
      -- CP-element group 12: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Update/cr
      -- 
    ra_10869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4394_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(12)); -- 
    cr_10873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(12), ack => RPIPE_Block7_starting_4394_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4394_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Sample/rr
      -- 
    ca_10874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4394_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(13)); -- 
    rr_10882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(13), ack => RPIPE_Block7_starting_4397_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_update_start_
      -- CP-element group 14: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Update/cr
      -- 
    ra_10883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4397_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(14)); -- 
    cr_10887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(14), ack => RPIPE_Block7_starting_4397_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	32 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	33 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15:  members (61) 
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/$exit
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398__exit__
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519__entry__
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4380_to_assign_stmt_4398/RPIPE_Block7_starting_4397_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_update_start_
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Update/cr
      -- 
    ca_10888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block7_starting_4397_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(15)); -- 
    rr_10899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4402_inst_req_0); -- 
    cr_10904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4402_inst_req_1); -- 
    rr_10913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4412_inst_req_0); -- 
    cr_10918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4412_inst_req_1); -- 
    rr_10927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4428_inst_req_0); -- 
    cr_10932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4428_inst_req_1); -- 
    rr_10941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4432_inst_req_0); -- 
    cr_10946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4432_inst_req_1); -- 
    rr_10955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4436_inst_req_0); -- 
    cr_10960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4436_inst_req_1); -- 
    rr_10969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4440_inst_req_0); -- 
    cr_10974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4440_inst_req_1); -- 
    rr_10983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4449_inst_req_0); -- 
    cr_10988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4449_inst_req_1); -- 
    rr_10997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4453_inst_req_0); -- 
    cr_11002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4453_inst_req_1); -- 
    rr_11011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4483_inst_req_0); -- 
    cr_11016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(15), ack => type_cast_4483_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Sample/ra
      -- 
    ra_10900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4402_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4402_Update/ca
      -- 
    ca_10905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4402_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Sample/ra
      -- 
    ra_10914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4412_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4412_Update/ca
      -- 
    ca_10919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4412_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Sample/ra
      -- 
    ra_10928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4428_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4428_Update/ca
      -- 
    ca_10933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4428_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Sample/ra
      -- 
    ra_10942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4432_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4432_Update/ca
      -- 
    ca_10947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4432_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Sample/ra
      -- 
    ra_10956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4436_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4436_Update/ca
      -- 
    ca_10961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4436_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Sample/ra
      -- 
    ra_10970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4440_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4440_Update/ca
      -- 
    ca_10975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4440_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Sample/ra
      -- 
    ra_10984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4449_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4449_Update/ca
      -- 
    ca_10989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4449_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Sample/ra
      -- 
    ra_10998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4453_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4453_Update/ca
      -- 
    ca_11003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4453_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Sample/ra
      -- 
    ra_11012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4483_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/type_cast_4483_Update/ca
      -- 
    ca_11017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4483_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	19 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	91 
    -- CP-element group 34: 	92 
    -- CP-element group 34: 	93 
    -- CP-element group 34: 	95 
    -- CP-element group 34: 	96 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519__exit__
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_4377/assign_stmt_4403_to_assign_stmt_4519/$exit
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4522/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Update/cr
      -- 
    rr_11614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(34), ack => type_cast_4532_inst_req_0); -- 
    cr_11619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(34), ack => type_cast_4532_inst_req_1); -- 
    rr_11637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(34), ack => type_cast_4538_inst_req_0); -- 
    cr_11642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(34), ack => type_cast_4538_inst_req_1); -- 
    zeropad3D_H_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(31) & zeropad3D_H_CP_10732_elements(33) & zeropad3D_H_CP_10732_elements(17) & zeropad3D_H_CP_10732_elements(19) & zeropad3D_H_CP_10732_elements(21) & zeropad3D_H_CP_10732_elements(23) & zeropad3D_H_CP_10732_elements(25) & zeropad3D_H_CP_10732_elements(27) & zeropad3D_H_CP_10732_elements(29);
      gj_zeropad3D_H_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	113 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Sample/ra
      -- 
    ra_11029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4545_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	113 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (13) 
      -- CP-element group 36: 	 branch_block_stmt_4377/R_orx_xcond_4573_place
      -- CP-element group 36: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571__exit__
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572__entry__
      -- CP-element group 36: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/$exit
      -- CP-element group 36: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_4377/if_stmt_4572_else_link/$entry
      -- 
    ca_11034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4545_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(36)); -- 
    branch_req_11042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(36), ack => if_stmt_4572_branch_req_0); -- 
    -- CP-element group 37:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	40 
    -- CP-element group 37:  members (18) 
      -- CP-element group 37: 	 branch_block_stmt_4377/whilex_xbody_lorx_xlhsx_xfalse64
      -- CP-element group 37: 	 branch_block_stmt_4377/merge_stmt_4578_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_4377/whilex_xbody_lorx_xlhsx_xfalse64_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_4377/whilex_xbody_lorx_xlhsx_xfalse64_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_4377/merge_stmt_4578_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_4377/merge_stmt_4578_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_4377/merge_stmt_4578__exit__
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608__entry__
      -- CP-element group 37: 	 branch_block_stmt_4377/if_stmt_4572_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_4377/if_stmt_4572_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/$entry
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_update_start_
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_4377/merge_stmt_4578_PhiAck/dummy
      -- 
    if_choice_transition_11047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4572_branch_ack_1, ack => zeropad3D_H_CP_10732_elements(37)); -- 
    rr_11064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(37), ack => type_cast_4582_inst_req_0); -- 
    cr_11069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(37), ack => type_cast_4582_inst_req_1); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	114 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_4377/whilex_xbody_ifx_xthen
      -- CP-element group 38: 	 branch_block_stmt_4377/if_stmt_4572_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_4377/if_stmt_4572_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_4377/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 38: 	 branch_block_stmt_4377/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- 
    else_choice_transition_11051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4572_branch_ack_0, ack => zeropad3D_H_CP_10732_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Sample/ra
      -- 
    ra_11065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4582_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(39)); -- 
    -- CP-element group 40:  branch  transition  place  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (13) 
      -- CP-element group 40: 	 branch_block_stmt_4377/R_orx_xcond193_4610_place
      -- CP-element group 40: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608__exit__
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609__entry__
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609_else_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/$exit
      -- CP-element group 40: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_4377/assign_stmt_4583_to_assign_stmt_4608/type_cast_4582_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609_dead_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609_eval_test/$entry
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609_eval_test/$exit
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609_eval_test/branch_req
      -- CP-element group 40: 	 branch_block_stmt_4377/if_stmt_4609_if_link/$entry
      -- 
    ca_11070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4582_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(40)); -- 
    branch_req_11078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(40), ack => if_stmt_4609_branch_req_0); -- 
    -- CP-element group 41:  fork  transition  place  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	64 
    -- CP-element group 41: 	62 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	58 
    -- CP-element group 41: 	60 
    -- CP-element group 41: 	66 
    -- CP-element group 41: 	68 
    -- CP-element group 41: 	70 
    -- CP-element group 41: 	72 
    -- CP-element group 41: 	75 
    -- CP-element group 41:  members (46) 
      -- CP-element group 41: 	 branch_block_stmt_4377/merge_stmt_4673_PhiReqMerge
      -- CP-element group 41: 	 branch_block_stmt_4377/merge_stmt_4673__exit__
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778__entry__
      -- CP-element group 41: 	 branch_block_stmt_4377/if_stmt_4609_if_link/$exit
      -- CP-element group 41: 	 branch_block_stmt_4377/if_stmt_4609_if_link/if_choice_transition
      -- CP-element group 41: 	 branch_block_stmt_4377/lorx_xlhsx_xfalse64_ifx_xelse
      -- CP-element group 41: 	 branch_block_stmt_4377/merge_stmt_4673_PhiAck/dummy
      -- CP-element group 41: 	 branch_block_stmt_4377/merge_stmt_4673_PhiAck/$exit
      -- CP-element group 41: 	 branch_block_stmt_4377/merge_stmt_4673_PhiAck/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/lorx_xlhsx_xfalse64_ifx_xelse_PhiReq/$exit
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/lorx_xlhsx_xfalse64_ifx_xelse_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_complete/req
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_complete/req
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_update_start_
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/word_access_complete/word_0/cr
      -- 
    if_choice_transition_11083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4609_branch_ack_1, ack => zeropad3D_H_CP_10732_elements(41)); -- 
    rr_11241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => type_cast_4677_inst_req_0); -- 
    cr_11246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => type_cast_4677_inst_req_1); -- 
    cr_11260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => type_cast_4741_inst_req_1); -- 
    req_11291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => array_obj_ref_4747_index_offset_req_1); -- 
    req_11306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => addr_of_4748_final_reg_req_1); -- 
    cr_11351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => ptr_deref_4752_load_0_req_1); -- 
    cr_11370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => type_cast_4766_inst_req_1); -- 
    req_11401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => array_obj_ref_4772_index_offset_req_1); -- 
    req_11416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => addr_of_4773_final_reg_req_1); -- 
    cr_11466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(41), ack => ptr_deref_4776_store_0_req_1); -- 
    -- CP-element group 42:  transition  place  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	114 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_4377/if_stmt_4609_else_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_4377/if_stmt_4609_else_link/else_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_4377/lorx_xlhsx_xfalse64_ifx_xthen
      -- CP-element group 42: 	 branch_block_stmt_4377/lorx_xlhsx_xfalse64_ifx_xthen_PhiReq/$exit
      -- CP-element group 42: 	 branch_block_stmt_4377/lorx_xlhsx_xfalse64_ifx_xthen_PhiReq/$entry
      -- 
    else_choice_transition_11087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4609_branch_ack_0, ack => zeropad3D_H_CP_10732_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	114 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Sample/ra
      -- 
    ra_11101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4619_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	114 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Update/ca
      -- 
    ca_11106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4619_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	114 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Sample/ra
      -- 
    ra_11115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4624_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	114 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Update/ca
      -- 
    ca_11120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4624_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Sample/rr
      -- 
    rr_11128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(47), ack => type_cast_4658_inst_req_0); -- 
    zeropad3D_H_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(46) & zeropad3D_H_CP_10732_elements(44);
      gj_zeropad3D_H_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Sample/ra
      -- 
    ra_11129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4658_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	114 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Sample/req
      -- 
    ca_11134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4658_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(49)); -- 
    req_11159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(49), ack => array_obj_ref_4664_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	56 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Sample/ack
      -- 
    ack_11160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4664_index_offset_ack_0, ack => zeropad3D_H_CP_10732_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	114 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_request/req
      -- 
    ack_11165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4664_index_offset_ack_1, ack => zeropad3D_H_CP_10732_elements(51)); -- 
    req_11174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(51), ack => addr_of_4665_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_request/ack
      -- 
    ack_11175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4665_final_reg_ack_0, ack => zeropad3D_H_CP_10732_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	114 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (28) 
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/ptr_deref_4668_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/ptr_deref_4668_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/ptr_deref_4668_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/ptr_deref_4668_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/word_access_start/word_0/rr
      -- 
    ack_11180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4665_final_reg_ack_1, ack => zeropad3D_H_CP_10732_elements(53)); -- 
    rr_11218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(53), ack => ptr_deref_4668_store_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Sample/word_access_start/word_0/ra
      -- 
    ra_11219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4668_store_0_ack_0, ack => zeropad3D_H_CP_10732_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	114 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/word_access_complete/word_0/ca
      -- 
    ca_11230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4668_store_0_ack_1, ack => zeropad3D_H_CP_10732_elements(55)); -- 
    -- CP-element group 56:  join  transition  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	50 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	115 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_4377/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_4377/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671__exit__
      -- CP-element group 56: 	 branch_block_stmt_4377/ifx_xthen_ifx_xend
      -- CP-element group 56: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/$exit
      -- 
    zeropad3D_H_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(50) & zeropad3D_H_CP_10732_elements(55);
      gj_zeropad3D_H_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Sample/ra
      -- 
    ra_11242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4677_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	67 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4677_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Sample/rr
      -- 
    ca_11247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4677_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(58)); -- 
    rr_11255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(58), ack => type_cast_4741_inst_req_0); -- 
    rr_11365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(58), ack => type_cast_4766_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Sample/ra
      -- 
    ra_11256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4741_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	41 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (16) 
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4741_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_scale_1/scale_rename_req
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Sample/req
      -- 
    ca_11261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4741_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(60)); -- 
    req_11286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(60), ack => array_obj_ref_4747_index_offset_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	76 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Sample/ack
      -- 
    ack_11287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4747_index_offset_ack_0, ack => zeropad3D_H_CP_10732_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	41 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (11) 
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_offset_calculated
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_final_index_sum_regn_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4747_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_request/$entry
      -- CP-element group 62: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_request/req
      -- 
    ack_11292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4747_index_offset_ack_1, ack => zeropad3D_H_CP_10732_elements(62)); -- 
    req_11301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(62), ack => addr_of_4748_final_reg_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_request/$exit
      -- CP-element group 63: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_request/ack
      -- 
    ack_11302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4748_final_reg_ack_0, ack => zeropad3D_H_CP_10732_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	41 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (24) 
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4748_complete/ack
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_word_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_address_resized
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_addr_resize/$entry
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_addr_resize/$exit
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_addr_resize/base_resize_req
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_addr_resize/base_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_word_addrgen/$entry
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_word_addrgen/$exit
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_word_addrgen/root_register_req
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_word_addrgen/root_register_ack
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/word_access_start/word_0/rr
      -- 
    ack_11307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4748_final_reg_ack_1, ack => zeropad3D_H_CP_10732_elements(64)); -- 
    rr_11340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(64), ack => ptr_deref_4752_load_0_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Sample/word_access_start/word_0/ra
      -- 
    ra_11341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4752_load_0_ack_0, ack => zeropad3D_H_CP_10732_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	41 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	73 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/word_access_complete/word_0/ca
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/ptr_deref_4752_Merge/$entry
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/ptr_deref_4752_Merge/$exit
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/ptr_deref_4752_Merge/merge_req
      -- CP-element group 66: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4752_Update/ptr_deref_4752_Merge/merge_ack
      -- 
    ca_11352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4752_load_0_ack_1, ack => zeropad3D_H_CP_10732_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	58 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Sample/ra
      -- 
    ra_11366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4766_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	41 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/type_cast_4766_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_resized_1
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_scaled_1
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_computed_1
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_resize_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_resize_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_resize_1/index_resize_req
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_resize_1/index_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_scale_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_scale_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_scale_1/scale_rename_req
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_index_scale_1/scale_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Sample/req
      -- 
    ca_11371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4766_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(68)); -- 
    req_11396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(68), ack => array_obj_ref_4772_index_offset_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	76 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_sample_complete
      -- CP-element group 69: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Sample/ack
      -- 
    ack_11397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4772_index_offset_ack_0, ack => zeropad3D_H_CP_10732_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	41 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (11) 
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_offset_calculated
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_final_index_sum_regn_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/array_obj_ref_4772_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_request/$entry
      -- CP-element group 70: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_request/req
      -- 
    ack_11402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4772_index_offset_ack_1, ack => zeropad3D_H_CP_10732_elements(70)); -- 
    req_11411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(70), ack => addr_of_4773_final_reg_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_request/$exit
      -- CP-element group 71: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_request/ack
      -- 
    ack_11412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4773_final_reg_ack_0, ack => zeropad3D_H_CP_10732_elements(71)); -- 
    -- CP-element group 72:  fork  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	41 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (19) 
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/addr_of_4773_complete/ack
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_word_addrgen/root_register_ack
      -- 
    ack_11417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4773_final_reg_ack_1, ack => zeropad3D_H_CP_10732_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/ptr_deref_4776_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/ptr_deref_4776_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/ptr_deref_4776_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/ptr_deref_4776_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/word_access_start/word_0/rr
      -- 
    rr_11455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(73), ack => ptr_deref_4776_store_0_req_0); -- 
    zeropad3D_H_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(66) & zeropad3D_H_CP_10732_elements(72);
      gj_zeropad3D_H_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Sample/word_access_start/word_0/ra
      -- 
    ra_11456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4776_store_0_ack_0, ack => zeropad3D_H_CP_10732_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/ptr_deref_4776_Update/word_access_complete/word_0/ca
      -- 
    ca_11467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4776_store_0_ack_1, ack => zeropad3D_H_CP_10732_elements(75)); -- 
    -- CP-element group 76:  join  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	61 
    -- CP-element group 76: 	69 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	115 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_4377/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_4377/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778__exit__
      -- CP-element group 76: 	 branch_block_stmt_4377/ifx_xelse_ifx_xend
      -- CP-element group 76: 	 branch_block_stmt_4377/assign_stmt_4678_to_assign_stmt_4778/$exit
      -- 
    zeropad3D_H_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(61) & zeropad3D_H_CP_10732_elements(69) & zeropad3D_H_CP_10732_elements(75);
      gj_zeropad3D_H_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	115 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Sample/ra
      -- 
    ra_11479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4784_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(77)); -- 
    -- CP-element group 78:  branch  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	115 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (13) 
      -- CP-element group 78: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798__exit__
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799__entry__
      -- CP-element group 78: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/$exit
      -- CP-element group 78: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799_dead_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799_eval_test/$entry
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799_eval_test/$exit
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799_eval_test/branch_req
      -- CP-element group 78: 	 branch_block_stmt_4377/R_cmp148_4800_place
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799_if_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_4377/if_stmt_4799_else_link/$entry
      -- 
    ca_11484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4784_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(78)); -- 
    branch_req_11492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(78), ack => if_stmt_4799_branch_req_0); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	124 
    -- CP-element group 79: 	125 
    -- CP-element group 79: 	127 
    -- CP-element group 79: 	128 
    -- CP-element group 79: 	130 
    -- CP-element group 79: 	131 
    -- CP-element group 79:  members (40) 
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xend_ifx_xthen150_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_4377/merge_stmt_4805_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xend_ifx_xthen150_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/merge_stmt_4805_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_4377/merge_stmt_4805_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/merge_stmt_4805__exit__
      -- CP-element group 79: 	 branch_block_stmt_4377/assign_stmt_4811__entry__
      -- CP-element group 79: 	 branch_block_stmt_4377/assign_stmt_4811__exit__
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/merge_stmt_4805_PhiAck/dummy
      -- CP-element group 79: 	 branch_block_stmt_4377/if_stmt_4799_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_4377/if_stmt_4799_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_4377/ifx_xend_ifx_xthen150
      -- CP-element group 79: 	 branch_block_stmt_4377/assign_stmt_4811/$entry
      -- CP-element group 79: 	 branch_block_stmt_4377/assign_stmt_4811/$exit
      -- 
    if_choice_transition_11497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4799_branch_ack_1, ack => zeropad3D_H_CP_10732_elements(79)); -- 
    cr_11920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(79), ack => type_cast_4868_inst_req_1); -- 
    rr_11869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(79), ack => type_cast_4878_inst_req_0); -- 
    rr_11915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(79), ack => type_cast_4868_inst_req_0); -- 
    rr_11892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(79), ack => type_cast_4872_inst_req_0); -- 
    cr_11874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(79), ack => type_cast_4878_inst_req_1); -- 
    cr_11897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(79), ack => type_cast_4872_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  place  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80: 	84 
    -- CP-element group 80: 	86 
    -- CP-element group 80:  members (24) 
      -- CP-element group 80: 	 branch_block_stmt_4377/merge_stmt_4813_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_4377/merge_stmt_4813__exit__
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854__entry__
      -- CP-element group 80: 	 branch_block_stmt_4377/merge_stmt_4813_PhiAck/dummy
      -- CP-element group 80: 	 branch_block_stmt_4377/merge_stmt_4813_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_4377/merge_stmt_4813_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/ifx_xend_ifx_xelse155_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_4377/ifx_xend_ifx_xelse155_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/if_stmt_4799_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_4377/if_stmt_4799_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_4377/ifx_xend_ifx_xelse155
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_update_start_
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_update_start_
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_update_start_
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Update/cr
      -- 
    else_choice_transition_11501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4799_branch_ack_0, ack => zeropad3D_H_CP_10732_elements(80)); -- 
    rr_11517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(80), ack => type_cast_4823_inst_req_0); -- 
    cr_11522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(80), ack => type_cast_4823_inst_req_1); -- 
    cr_11536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(80), ack => type_cast_4832_inst_req_1); -- 
    cr_11550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(80), ack => type_cast_4848_inst_req_1); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Sample/ra
      -- 
    ra_11518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4823_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4823_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Sample/rr
      -- 
    ca_11523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4823_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(82)); -- 
    rr_11531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(82), ack => type_cast_4832_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Sample/ra
      -- 
    ra_11532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4832_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4832_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Sample/rr
      -- 
    ca_11537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4832_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(84)); -- 
    rr_11545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(84), ack => type_cast_4848_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Sample/ra
      -- 
    ra_11546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4848_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(85)); -- 
    -- CP-element group 86:  branch  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	80 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (13) 
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855__entry__
      -- CP-element group 86: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854__exit__
      -- CP-element group 86: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/$exit
      -- CP-element group 86: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_4377/assign_stmt_4819_to_assign_stmt_4854/type_cast_4848_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_4377/R_cmp179_4856_place
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_4377/if_stmt_4855_else_link/$entry
      -- 
    ca_11551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4848_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(86)); -- 
    branch_req_11559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(86), ack => if_stmt_4855_branch_req_0); -- 
    -- CP-element group 87:  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (15) 
      -- CP-element group 87: 	 branch_block_stmt_4377/assign_stmt_4888__entry__
      -- CP-element group 87: 	 branch_block_stmt_4377/merge_stmt_4883__exit__
      -- CP-element group 87: 	 branch_block_stmt_4377/merge_stmt_4883_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_4377/merge_stmt_4883_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_4377/merge_stmt_4883_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_4377/merge_stmt_4883_PhiAck/dummy
      -- CP-element group 87: 	 branch_block_stmt_4377/ifx_xelse155_whilex_xend_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_4377/ifx_xelse155_whilex_xend_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_4377/if_stmt_4855_if_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_4377/if_stmt_4855_if_link/if_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_4377/ifx_xelse155_whilex_xend
      -- CP-element group 87: 	 branch_block_stmt_4377/assign_stmt_4888/$entry
      -- CP-element group 87: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Sample/req
      -- 
    if_choice_transition_11564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4855_branch_ack_1, ack => zeropad3D_H_CP_10732_elements(87)); -- 
    req_11581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(87), ack => WPIPE_Block7_complete_4885_inst_req_0); -- 
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	116 
    -- CP-element group 88: 	117 
    -- CP-element group 88: 	119 
    -- CP-element group 88: 	120 
    -- CP-element group 88: 	122 
    -- CP-element group 88:  members (22) 
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4862/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_4377/if_stmt_4855_else_link/$exit
      -- CP-element group 88: 	 branch_block_stmt_4377/if_stmt_4855_else_link/else_choice_transition
      -- CP-element group 88: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187
      -- 
    else_choice_transition_11568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4855_branch_ack_0, ack => zeropad3D_H_CP_10732_elements(88)); -- 
    rr_11835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(88), ack => type_cast_4874_inst_req_0); -- 
    rr_11812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(88), ack => type_cast_4880_inst_req_0); -- 
    cr_11840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(88), ack => type_cast_4874_inst_req_1); -- 
    cr_11817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(88), ack => type_cast_4880_inst_req_1); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_update_start_
      -- CP-element group 89: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Update/req
      -- 
    ack_11582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_complete_4885_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(89)); -- 
    req_11586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(89), ack => WPIPE_Block7_complete_4885_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (16) 
      -- CP-element group 90: 	 branch_block_stmt_4377/merge_stmt_4890__exit__
      -- CP-element group 90: 	 branch_block_stmt_4377/return__
      -- CP-element group 90: 	 branch_block_stmt_4377/assign_stmt_4888__exit__
      -- CP-element group 90: 	 branch_block_stmt_4377/merge_stmt_4890_PhiAck/dummy
      -- CP-element group 90: 	 branch_block_stmt_4377/merge_stmt_4890_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_4377/merge_stmt_4890_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_4377/merge_stmt_4890_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_4377/return___PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_4377/return___PhiReq/$exit
      -- CP-element group 90: 	 $exit
      -- CP-element group 90: 	 branch_block_stmt_4377/$exit
      -- CP-element group 90: 	 branch_block_stmt_4377/branch_block_stmt_4377__exit__
      -- CP-element group 90: 	 branch_block_stmt_4377/assign_stmt_4888/$exit
      -- CP-element group 90: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_4377/assign_stmt_4888/WPIPE_Block7_complete_4885_Update/ack
      -- 
    ack_11587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block7_complete_4885_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(90)); -- 
    -- CP-element group 91:  transition  output  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	34 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4522/$exit
      -- CP-element group 91: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4526_konst_delay_trans
      -- CP-element group 91: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_req
      -- 
    phi_stmt_4522_req_11598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4522_req_11598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(91), ack => phi_stmt_4522_req_0); -- 
    -- Element group zeropad3D_H_CP_10732_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => zeropad3D_H_CP_10732_elements(34), ack => zeropad3D_H_CP_10732_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	34 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Sample/ra
      -- 
    ra_11615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4532_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	34 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/Update/ca
      -- 
    ca_11620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4532_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/$exit
      -- CP-element group 94: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/$exit
      -- CP-element group 94: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4532/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_req
      -- 
    phi_stmt_4529_req_11621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4529_req_11621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(94), ack => phi_stmt_4529_req_0); -- 
    zeropad3D_H_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(92) & zeropad3D_H_CP_10732_elements(93);
      gj_zeropad3D_H_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	34 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Sample/ra
      -- 
    ra_11638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4538_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	34 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/Update/ca
      -- 
    ca_11643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4538_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/$exit
      -- CP-element group 97: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/$exit
      -- CP-element group 97: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4538/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_req
      -- 
    phi_stmt_4535_req_11644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4535_req_11644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(97), ack => phi_stmt_4535_req_0); -- 
    zeropad3D_H_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(95) & zeropad3D_H_CP_10732_elements(96);
      gj_zeropad3D_H_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	109 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_4377/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_H_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_H_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(91) & zeropad3D_H_CP_10732_elements(94) & zeropad3D_H_CP_10732_elements(97);
      gj_zeropad3D_H_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Sample/$exit
      -- 
    ra_11664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4528_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Update/ca
      -- CP-element group 100: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/Update/$exit
      -- 
    ca_11669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4528_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_req
      -- CP-element group 101: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/$exit
      -- CP-element group 101: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/$exit
      -- CP-element group 101: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4522/phi_stmt_4522_sources/type_cast_4528/SplitProtocol/$exit
      -- 
    phi_stmt_4522_req_11670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4522_req_11670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(101), ack => phi_stmt_4522_req_1); -- 
    zeropad3D_H_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(99) & zeropad3D_H_CP_10732_elements(100);
      gj_zeropad3D_H_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Sample/ra
      -- 
    ra_11687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4534_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/Update/ca
      -- 
    ca_11692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4534_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/$exit
      -- CP-element group 104: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_req
      -- CP-element group 104: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/$exit
      -- CP-element group 104: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4529/phi_stmt_4529_sources/type_cast_4534/SplitProtocol/$exit
      -- 
    phi_stmt_4529_req_11693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4529_req_11693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(104), ack => phi_stmt_4529_req_1); -- 
    zeropad3D_H_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(102) & zeropad3D_H_CP_10732_elements(103);
      gj_zeropad3D_H_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	1 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Sample/ra
      -- 
    ra_11710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4540_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/Update/ca
      -- 
    ca_11715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4540_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_req
      -- CP-element group 107: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/$exit
      -- CP-element group 107: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/type_cast_4540/$exit
      -- CP-element group 107: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/phi_stmt_4535/phi_stmt_4535_sources/$exit
      -- 
    phi_stmt_4535_req_11716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4535_req_11716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(107), ack => phi_stmt_4535_req_1); -- 
    zeropad3D_H_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(105) & zeropad3D_H_CP_10732_elements(106);
      gj_zeropad3D_H_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_4377/ifx_xend187_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_H_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(101) & zeropad3D_H_CP_10732_elements(104) & zeropad3D_H_CP_10732_elements(107);
      gj_zeropad3D_H_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	98 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_4377/merge_stmt_4521_PhiAck/$entry
      -- CP-element group 109: 	 branch_block_stmt_4377/merge_stmt_4521_PhiReqMerge
      -- 
    zeropad3D_H_CP_10732_elements(109) <= OrReduce(zeropad3D_H_CP_10732_elements(98) & zeropad3D_H_CP_10732_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_4377/merge_stmt_4521_PhiAck/phi_stmt_4522_ack
      -- 
    phi_stmt_4522_ack_11721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4522_ack_0, ack => zeropad3D_H_CP_10732_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_4377/merge_stmt_4521_PhiAck/phi_stmt_4529_ack
      -- 
    phi_stmt_4529_ack_11722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4529_ack_0, ack => zeropad3D_H_CP_10732_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_4377/merge_stmt_4521_PhiAck/phi_stmt_4535_ack
      -- 
    phi_stmt_4535_ack_11723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4535_ack_0, ack => zeropad3D_H_CP_10732_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	35 
    -- CP-element group 113: 	36 
    -- CP-element group 113:  members (10) 
      -- CP-element group 113: 	 branch_block_stmt_4377/merge_stmt_4521_PhiAck/$exit
      -- CP-element group 113: 	 branch_block_stmt_4377/merge_stmt_4521__exit__
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571__entry__
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/$entry
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_update_start_
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_4377/assign_stmt_4546_to_assign_stmt_4571/type_cast_4545_Update/cr
      -- 
    rr_11028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(113), ack => type_cast_4545_inst_req_0); -- 
    cr_11033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(113), ack => type_cast_4545_inst_req_1); -- 
    zeropad3D_H_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(110) & zeropad3D_H_CP_10732_elements(111) & zeropad3D_H_CP_10732_elements(112);
      gj_zeropad3D_H_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  merge  fork  transition  place  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	38 
    -- CP-element group 114: 	42 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	51 
    -- CP-element group 114: 	53 
    -- CP-element group 114: 	45 
    -- CP-element group 114: 	46 
    -- CP-element group 114: 	55 
    -- CP-element group 114: 	49 
    -- CP-element group 114: 	43 
    -- CP-element group 114: 	44 
    -- CP-element group 114:  members (33) 
      -- CP-element group 114: 	 branch_block_stmt_4377/merge_stmt_4615_PhiReqMerge
      -- CP-element group 114: 	 branch_block_stmt_4377/merge_stmt_4615__exit__
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671__entry__
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_update_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4619_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_update_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4624_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_update_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/type_cast_4658_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_update_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_update_start
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/array_obj_ref_4664_final_index_sum_regn_Update/req
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/addr_of_4665_complete/req
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_update_start_
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/word_access_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/word_access_complete/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_4377/assign_stmt_4620_to_assign_stmt_4671/ptr_deref_4668_Update/word_access_complete/word_0/cr
      -- CP-element group 114: 	 branch_block_stmt_4377/merge_stmt_4615_PhiAck/dummy
      -- CP-element group 114: 	 branch_block_stmt_4377/merge_stmt_4615_PhiAck/$exit
      -- CP-element group 114: 	 branch_block_stmt_4377/merge_stmt_4615_PhiAck/$entry
      -- 
    rr_11100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => type_cast_4619_inst_req_0); -- 
    cr_11105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => type_cast_4619_inst_req_1); -- 
    rr_11114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => type_cast_4624_inst_req_0); -- 
    cr_11119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => type_cast_4624_inst_req_1); -- 
    cr_11133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => type_cast_4658_inst_req_1); -- 
    req_11164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => array_obj_ref_4664_index_offset_req_1); -- 
    req_11179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => addr_of_4665_final_reg_req_1); -- 
    cr_11229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(114), ack => ptr_deref_4668_store_0_req_1); -- 
    zeropad3D_H_CP_10732_elements(114) <= OrReduce(zeropad3D_H_CP_10732_elements(38) & zeropad3D_H_CP_10732_elements(42));
    -- CP-element group 115:  merge  fork  transition  place  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	56 
    -- CP-element group 115: 	76 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	77 
    -- CP-element group 115: 	78 
    -- CP-element group 115:  members (13) 
      -- CP-element group 115: 	 branch_block_stmt_4377/merge_stmt_4780_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_4377/merge_stmt_4780_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_4377/merge_stmt_4780_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_4377/merge_stmt_4780_PhiAck/dummy
      -- CP-element group 115: 	 branch_block_stmt_4377/merge_stmt_4780__exit__
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798__entry__
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/$entry
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_update_start_
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_4377/assign_stmt_4785_to_assign_stmt_4798/type_cast_4784_Update/cr
      -- 
    rr_11478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(115), ack => type_cast_4784_inst_req_0); -- 
    cr_11483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(115), ack => type_cast_4784_inst_req_1); -- 
    zeropad3D_H_CP_10732_elements(115) <= OrReduce(zeropad3D_H_CP_10732_elements(56) & zeropad3D_H_CP_10732_elements(76));
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	88 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Sample/ra
      -- 
    ra_11813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4880_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	88 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/Update/ca
      -- 
    ca_11818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4880_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/$exit
      -- CP-element group 118: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/$exit
      -- CP-element group 118: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4880/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_req
      -- 
    phi_stmt_4875_req_11819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4875_req_11819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(118), ack => phi_stmt_4875_req_1); -- 
    zeropad3D_H_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(116) & zeropad3D_H_CP_10732_elements(117);
      gj_zeropad3D_H_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	88 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Sample/ra
      -- 
    ra_11836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4874_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	88 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/Update/ca
      -- 
    ca_11841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4874_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4874/$exit
      -- CP-element group 121: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_req
      -- CP-element group 121: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4869/$exit
      -- 
    phi_stmt_4869_req_11842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4869_req_11842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(121), ack => phi_stmt_4869_req_1); -- 
    zeropad3D_H_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(119) & zeropad3D_H_CP_10732_elements(120);
      gj_zeropad3D_H_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  output  delay-element  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	88 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4862/$exit
      -- CP-element group 122: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_req
      -- CP-element group 122: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4866_konst_delay_trans
      -- CP-element group 122: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/$exit
      -- 
    phi_stmt_4862_req_11850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4862_req_11850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(122), ack => phi_stmt_4862_req_0); -- 
    -- Element group zeropad3D_H_CP_10732_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => zeropad3D_H_CP_10732_elements(88), ack => zeropad3D_H_CP_10732_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	134 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_4377/ifx_xelse155_ifx_xend187_PhiReq/$exit
      -- 
    zeropad3D_H_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(118) & zeropad3D_H_CP_10732_elements(121) & zeropad3D_H_CP_10732_elements(122);
      gj_zeropad3D_H_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	79 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Sample/ra
      -- 
    ra_11870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4878_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/Update/ca
      -- 
    ca_11875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4878_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	133 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/SplitProtocol/$exit
      -- CP-element group 126: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/$exit
      -- CP-element group 126: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_req
      -- CP-element group 126: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4875/phi_stmt_4875_sources/type_cast_4878/$exit
      -- 
    phi_stmt_4875_req_11876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4875_req_11876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(126), ack => phi_stmt_4875_req_0); -- 
    zeropad3D_H_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(124) & zeropad3D_H_CP_10732_elements(125);
      gj_zeropad3D_H_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	79 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Sample/ra
      -- 
    ra_11893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4872_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	79 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/Update/ca
      -- 
    ca_11898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4872_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/type_cast_4872/$exit
      -- CP-element group 129: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_req
      -- CP-element group 129: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/$exit
      -- CP-element group 129: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4869/phi_stmt_4869_sources/$exit
      -- 
    phi_stmt_4869_req_11899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4869_req_11899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(129), ack => phi_stmt_4869_req_0); -- 
    zeropad3D_H_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(127) & zeropad3D_H_CP_10732_elements(128);
      gj_zeropad3D_H_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	79 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Sample/ra
      -- 
    ra_11916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4868_inst_ack_0, ack => zeropad3D_H_CP_10732_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	79 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/Update/ca
      -- 
    ca_11921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4868_inst_ack_1, ack => zeropad3D_H_CP_10732_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/$exit
      -- CP-element group 132: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/type_cast_4868/SplitProtocol/$exit
      -- CP-element group 132: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/$exit
      -- CP-element group 132: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_sources/$exit
      -- CP-element group 132: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/phi_stmt_4862/phi_stmt_4862_req
      -- 
    phi_stmt_4862_req_11922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4862_req_11922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_H_CP_10732_elements(132), ack => phi_stmt_4862_req_1); -- 
    zeropad3D_H_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(130) & zeropad3D_H_CP_10732_elements(131);
      gj_zeropad3D_H_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	126 
    -- CP-element group 133: 	129 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_4377/ifx_xthen150_ifx_xend187_PhiReq/$exit
      -- 
    zeropad3D_H_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(126) & zeropad3D_H_CP_10732_elements(129) & zeropad3D_H_CP_10732_elements(132);
      gj_zeropad3D_H_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  merge  fork  transition  place  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	123 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_4377/merge_stmt_4861_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_4377/merge_stmt_4861_PhiAck/$entry
      -- 
    zeropad3D_H_CP_10732_elements(134) <= OrReduce(zeropad3D_H_CP_10732_elements(123) & zeropad3D_H_CP_10732_elements(133));
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_4377/merge_stmt_4861_PhiAck/phi_stmt_4862_ack
      -- 
    phi_stmt_4862_ack_11927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4862_ack_0, ack => zeropad3D_H_CP_10732_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_4377/merge_stmt_4861_PhiAck/phi_stmt_4869_ack
      -- 
    phi_stmt_4869_ack_11928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4869_ack_0, ack => zeropad3D_H_CP_10732_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_4377/merge_stmt_4861_PhiAck/phi_stmt_4875_ack
      -- 
    phi_stmt_4875_ack_11929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4875_ack_0, ack => zeropad3D_H_CP_10732_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	1 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_4377/merge_stmt_4861_PhiAck/$exit
      -- 
    zeropad3D_H_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_H_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_H_CP_10732_elements(135) & zeropad3D_H_CP_10732_elements(136) & zeropad3D_H_CP_10732_elements(137);
      gj_zeropad3D_H_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_H_CP_10732_elements(138), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_4467_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4517_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4652_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4735_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4760_wire : std_logic_vector(31 downto 0);
    signal R_idxprom135_4746_resized : std_logic_vector(13 downto 0);
    signal R_idxprom135_4746_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom140_4771_resized : std_logic_vector(13 downto 0);
    signal R_idxprom140_4771_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_4663_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_4663_scaled : std_logic_vector(13 downto 0);
    signal add107_4703 : std_logic_vector(31 downto 0);
    signal add116_4708 : std_logic_vector(31 downto 0);
    signal add126_4723 : std_logic_vector(31 downto 0);
    signal add132_4728 : std_logic_vector(31 downto 0);
    signal add145_4791 : std_logic_vector(31 downto 0);
    signal add153_4811 : std_logic_vector(15 downto 0);
    signal add163_4480 : std_logic_vector(31 downto 0);
    signal add178_4489 : std_logic_vector(31 downto 0);
    signal add78_4499 : std_logic_vector(31 downto 0);
    signal add89_4640 : std_logic_vector(31 downto 0);
    signal add95_4645 : std_logic_vector(31 downto 0);
    signal add_4494 : std_logic_vector(31 downto 0);
    signal array_obj_ref_4664_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4664_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4664_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4664_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4664_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4664_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4747_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4747_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4747_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4747_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4747_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4747_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4772_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4772_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4772_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4772_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4772_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4772_root_address : std_logic_vector(13 downto 0);
    signal arrayidx136_4749 : std_logic_vector(31 downto 0);
    signal arrayidx141_4774 : std_logic_vector(31 downto 0);
    signal arrayidx_4666 : std_logic_vector(31 downto 0);
    signal call1_4383 : std_logic_vector(7 downto 0);
    signal call2_4386 : std_logic_vector(7 downto 0);
    signal call3_4389 : std_logic_vector(7 downto 0);
    signal call4_4392 : std_logic_vector(7 downto 0);
    signal call5_4395 : std_logic_vector(7 downto 0);
    signal call6_4398 : std_logic_vector(7 downto 0);
    signal call_4380 : std_logic_vector(7 downto 0);
    signal cmp148_4798 : std_logic_vector(0 downto 0);
    signal cmp164_4829 : std_logic_vector(0 downto 0);
    signal cmp179_4854 : std_logic_vector(0 downto 0);
    signal cmp62_4566 : std_logic_vector(0 downto 0);
    signal cmp69_4590 : std_logic_vector(0 downto 0);
    signal cmp69x_xnot_4596 : std_logic_vector(0 downto 0);
    signal cmp79_4603 : std_logic_vector(0 downto 0);
    signal cmp_4553 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_4559 : std_logic_vector(0 downto 0);
    signal conv109_4519 : std_logic_vector(31 downto 0);
    signal conv10_4413 : std_logic_vector(15 downto 0);
    signal conv144_4785 : std_logic_vector(31 downto 0);
    signal conv158_4824 : std_logic_vector(31 downto 0);
    signal conv172_4849 : std_logic_vector(31 downto 0);
    signal conv174_4484 : std_logic_vector(31 downto 0);
    signal conv36_4429 : std_logic_vector(31 downto 0);
    signal conv38_4433 : std_logic_vector(31 downto 0);
    signal conv43_4437 : std_logic_vector(31 downto 0);
    signal conv45_4441 : std_logic_vector(31 downto 0);
    signal conv52_4546 : std_logic_vector(31 downto 0);
    signal conv54_4450 : std_logic_vector(31 downto 0);
    signal conv66_4583 : std_logic_vector(31 downto 0);
    signal conv83_4620 : std_logic_vector(31 downto 0);
    signal conv85_4454 : std_logic_vector(31 downto 0);
    signal conv87_4625 : std_logic_vector(31 downto 0);
    signal conv91_4469 : std_logic_vector(31 downto 0);
    signal conv99_4678 : std_logic_vector(31 downto 0);
    signal conv_4403 : std_logic_vector(15 downto 0);
    signal div11_4425 : std_logic_vector(15 downto 0);
    signal div_4409 : std_logic_vector(15 downto 0);
    signal idxprom135_4742 : std_logic_vector(63 downto 0);
    signal idxprom140_4767 : std_logic_vector(63 downto 0);
    signal idxprom_4659 : std_logic_vector(63 downto 0);
    signal inc169_4833 : std_logic_vector(15 downto 0);
    signal inc169x_xix_x2_4838 : std_logic_vector(15 downto 0);
    signal inc_4819 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_4869 : std_logic_vector(15 downto 0);
    signal ix_x2_4529 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_4875 : std_logic_vector(15 downto 0);
    signal jx_x1_4535 : std_logic_vector(15 downto 0);
    signal jx_x2_4844 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_4862 : std_logic_vector(15 downto 0);
    signal kx_x1_4522 : std_logic_vector(15 downto 0);
    signal mul106_4688 : std_logic_vector(31 downto 0);
    signal mul115_4698 : std_logic_vector(31 downto 0);
    signal mul125_4713 : std_logic_vector(31 downto 0);
    signal mul131_4718 : std_logic_vector(31 downto 0);
    signal mul39_4505 : std_logic_vector(31 downto 0);
    signal mul46_4446 : std_logic_vector(31 downto 0);
    signal mul88_4630 : std_logic_vector(31 downto 0);
    signal mul94_4635 : std_logic_vector(31 downto 0);
    signal mul_4419 : std_logic_vector(15 downto 0);
    signal orx_xcond193_4608 : std_logic_vector(0 downto 0);
    signal orx_xcond_4571 : std_logic_vector(0 downto 0);
    signal ptr_deref_4668_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4668_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4668_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4668_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4668_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4668_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4752_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4752_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4752_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4752_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4752_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4776_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4776_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4776_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4776_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4776_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4776_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext192_4460 : std_logic_vector(31 downto 0);
    signal sext_4510 : std_logic_vector(31 downto 0);
    signal shl_4475 : std_logic_vector(31 downto 0);
    signal shr134_4737 : std_logic_vector(31 downto 0);
    signal shr139_4762 : std_logic_vector(31 downto 0);
    signal shr_4654 : std_logic_vector(31 downto 0);
    signal sub114_4693 : std_logic_vector(31 downto 0);
    signal sub_4683 : std_logic_vector(31 downto 0);
    signal tmp137_4753 : std_logic_vector(63 downto 0);
    signal type_cast_4407_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4417_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4423_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4458_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4463_wire : std_logic_vector(31 downto 0);
    signal type_cast_4466_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4473_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4503_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4513_wire : std_logic_vector(31 downto 0);
    signal type_cast_4516_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4526_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4528_wire : std_logic_vector(15 downto 0);
    signal type_cast_4532_wire : std_logic_vector(15 downto 0);
    signal type_cast_4534_wire : std_logic_vector(15 downto 0);
    signal type_cast_4538_wire : std_logic_vector(15 downto 0);
    signal type_cast_4540_wire : std_logic_vector(15 downto 0);
    signal type_cast_4544_wire : std_logic_vector(31 downto 0);
    signal type_cast_4549_wire : std_logic_vector(31 downto 0);
    signal type_cast_4551_wire : std_logic_vector(31 downto 0);
    signal type_cast_4557_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_4562_wire : std_logic_vector(31 downto 0);
    signal type_cast_4564_wire : std_logic_vector(31 downto 0);
    signal type_cast_4581_wire : std_logic_vector(31 downto 0);
    signal type_cast_4586_wire : std_logic_vector(31 downto 0);
    signal type_cast_4588_wire : std_logic_vector(31 downto 0);
    signal type_cast_4594_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_4599_wire : std_logic_vector(31 downto 0);
    signal type_cast_4601_wire : std_logic_vector(31 downto 0);
    signal type_cast_4618_wire : std_logic_vector(31 downto 0);
    signal type_cast_4623_wire : std_logic_vector(31 downto 0);
    signal type_cast_4648_wire : std_logic_vector(31 downto 0);
    signal type_cast_4651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4657_wire : std_logic_vector(63 downto 0);
    signal type_cast_4670_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_4676_wire : std_logic_vector(31 downto 0);
    signal type_cast_4731_wire : std_logic_vector(31 downto 0);
    signal type_cast_4734_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4740_wire : std_logic_vector(63 downto 0);
    signal type_cast_4756_wire : std_logic_vector(31 downto 0);
    signal type_cast_4759_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4765_wire : std_logic_vector(63 downto 0);
    signal type_cast_4783_wire : std_logic_vector(31 downto 0);
    signal type_cast_4789_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4794_wire : std_logic_vector(31 downto 0);
    signal type_cast_4796_wire : std_logic_vector(31 downto 0);
    signal type_cast_4809_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4817_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4822_wire : std_logic_vector(31 downto 0);
    signal type_cast_4847_wire : std_logic_vector(31 downto 0);
    signal type_cast_4866_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4868_wire : std_logic_vector(15 downto 0);
    signal type_cast_4872_wire : std_logic_vector(15 downto 0);
    signal type_cast_4874_wire : std_logic_vector(15 downto 0);
    signal type_cast_4878_wire : std_logic_vector(15 downto 0);
    signal type_cast_4880_wire : std_logic_vector(15 downto 0);
    signal type_cast_4887_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_4664_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4664_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4664_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4664_resized_base_address <= "00000000000000";
    array_obj_ref_4747_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4747_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4747_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4747_resized_base_address <= "00000000000000";
    array_obj_ref_4772_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4772_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4772_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4772_resized_base_address <= "00000000000000";
    ptr_deref_4668_word_offset_0 <= "00000000000000";
    ptr_deref_4752_word_offset_0 <= "00000000000000";
    ptr_deref_4776_word_offset_0 <= "00000000000000";
    type_cast_4407_wire_constant <= "0000000000000001";
    type_cast_4417_wire_constant <= "0000000000000011";
    type_cast_4423_wire_constant <= "0000000000000010";
    type_cast_4458_wire_constant <= "00000000000000000000000000010000";
    type_cast_4466_wire_constant <= "00000000000000000000000000010000";
    type_cast_4473_wire_constant <= "00000000000000000000000000000001";
    type_cast_4503_wire_constant <= "00000000000000000000000000010000";
    type_cast_4516_wire_constant <= "00000000000000000000000000010000";
    type_cast_4526_wire_constant <= "0000000000000000";
    type_cast_4557_wire_constant <= "1";
    type_cast_4594_wire_constant <= "1";
    type_cast_4651_wire_constant <= "00000000000000000000000000000010";
    type_cast_4670_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4734_wire_constant <= "00000000000000000000000000000010";
    type_cast_4759_wire_constant <= "00000000000000000000000000000010";
    type_cast_4789_wire_constant <= "00000000000000000000000000000100";
    type_cast_4809_wire_constant <= "0000000000000100";
    type_cast_4817_wire_constant <= "0000000000000001";
    type_cast_4866_wire_constant <= "0000000000000000";
    type_cast_4887_wire_constant <= "00000001";
    phi_stmt_4522: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4526_wire_constant & type_cast_4528_wire;
      req <= phi_stmt_4522_req_0 & phi_stmt_4522_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4522",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4522_ack_0,
          idata => idata,
          odata => kx_x1_4522,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4522
    phi_stmt_4529: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4532_wire & type_cast_4534_wire;
      req <= phi_stmt_4529_req_0 & phi_stmt_4529_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4529",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4529_ack_0,
          idata => idata,
          odata => ix_x2_4529,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4529
    phi_stmt_4535: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4538_wire & type_cast_4540_wire;
      req <= phi_stmt_4535_req_0 & phi_stmt_4535_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4535",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4535_ack_0,
          idata => idata,
          odata => jx_x1_4535,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4535
    phi_stmt_4862: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4866_wire_constant & type_cast_4868_wire;
      req <= phi_stmt_4862_req_0 & phi_stmt_4862_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4862",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4862_ack_0,
          idata => idata,
          odata => kx_x0x_xph_4862,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4862
    phi_stmt_4869: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4872_wire & type_cast_4874_wire;
      req <= phi_stmt_4869_req_0 & phi_stmt_4869_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4869",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4869_ack_0,
          idata => idata,
          odata => ix_x1x_xph_4869,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4869
    phi_stmt_4875: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4878_wire & type_cast_4880_wire;
      req <= phi_stmt_4875_req_0 & phi_stmt_4875_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4875",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4875_ack_0,
          idata => idata,
          odata => jx_x0x_xph_4875,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4875
    -- flow-through select operator MUX_4843_inst
    jx_x2_4844 <= div_4409 when (cmp164_4829(0) /=  '0') else inc_4819;
    addr_of_4665_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4665_final_reg_req_0;
      addr_of_4665_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4665_final_reg_req_1;
      addr_of_4665_final_reg_ack_1<= rack(0);
      addr_of_4665_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4665_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4664_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_4666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4748_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4748_final_reg_req_0;
      addr_of_4748_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4748_final_reg_req_1;
      addr_of_4748_final_reg_ack_1<= rack(0);
      addr_of_4748_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4748_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4747_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx136_4749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4773_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4773_final_reg_req_0;
      addr_of_4773_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4773_final_reg_req_1;
      addr_of_4773_final_reg_ack_1<= rack(0);
      addr_of_4773_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4773_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4772_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx141_4774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4402_inst_req_0;
      type_cast_4402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4402_inst_req_1;
      type_cast_4402_inst_ack_1<= rack(0);
      type_cast_4402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_4383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_4403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4412_inst_req_0;
      type_cast_4412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4412_inst_req_1;
      type_cast_4412_inst_ack_1<= rack(0);
      type_cast_4412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_4380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_4413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4428_inst_req_0;
      type_cast_4428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4428_inst_req_1;
      type_cast_4428_inst_ack_1<= rack(0);
      type_cast_4428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_4386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_4429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4432_inst_req_0;
      type_cast_4432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4432_inst_req_1;
      type_cast_4432_inst_ack_1<= rack(0);
      type_cast_4432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_4383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_4433,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4436_inst_req_0;
      type_cast_4436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4436_inst_req_1;
      type_cast_4436_inst_ack_1<= rack(0);
      type_cast_4436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_4395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_4437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4440_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4440_inst_req_0;
      type_cast_4440_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4440_inst_req_1;
      type_cast_4440_inst_ack_1<= rack(0);
      type_cast_4440_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4440_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_4392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_4441,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4449_inst_req_0;
      type_cast_4449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4449_inst_req_1;
      type_cast_4449_inst_ack_1<= rack(0);
      type_cast_4449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_4398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_4450,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4453_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4453_inst_req_0;
      type_cast_4453_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4453_inst_req_1;
      type_cast_4453_inst_ack_1<= rack(0);
      type_cast_4453_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4453_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_4395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_4454,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4463_inst
    process(sext192_4460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext192_4460(31 downto 0);
      type_cast_4463_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4468_inst
    process(ASHR_i32_i32_4467_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4467_wire(31 downto 0);
      conv91_4469 <= tmp_var; -- 
    end process;
    type_cast_4483_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4483_inst_req_0;
      type_cast_4483_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4483_inst_req_1;
      type_cast_4483_inst_ack_1<= rack(0);
      type_cast_4483_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4483_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_4380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv174_4484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4513_inst
    process(sext_4510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_4510(31 downto 0);
      type_cast_4513_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4518_inst
    process(ASHR_i32_i32_4517_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4517_wire(31 downto 0);
      conv109_4519 <= tmp_var; -- 
    end process;
    type_cast_4528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4528_inst_req_0;
      type_cast_4528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4528_inst_req_1;
      type_cast_4528_inst_ack_1<= rack(0);
      type_cast_4528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_4862,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4528_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4532_inst_req_0;
      type_cast_4532_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4532_inst_req_1;
      type_cast_4532_inst_ack_1<= rack(0);
      type_cast_4532_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4532_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div11_4425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4532_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4534_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4534_inst_req_0;
      type_cast_4534_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4534_inst_req_1;
      type_cast_4534_inst_ack_1<= rack(0);
      type_cast_4534_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4534_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_4869,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4534_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4538_inst_req_0;
      type_cast_4538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4538_inst_req_1;
      type_cast_4538_inst_ack_1<= rack(0);
      type_cast_4538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_4409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4538_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4540_inst_req_0;
      type_cast_4540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4540_inst_req_1;
      type_cast_4540_inst_ack_1<= rack(0);
      type_cast_4540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_4875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4540_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4545_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4545_inst_req_0;
      type_cast_4545_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4545_inst_req_1;
      type_cast_4545_inst_ack_1<= rack(0);
      type_cast_4545_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4545_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4544_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_4546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4549_inst
    process(conv52_4546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv52_4546(31 downto 0);
      type_cast_4549_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4551_inst
    process(conv54_4450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv54_4450(31 downto 0);
      type_cast_4551_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4562_inst
    process(conv52_4546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv52_4546(31 downto 0);
      type_cast_4562_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4564_inst
    process(add_4494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_4494(31 downto 0);
      type_cast_4564_wire <= tmp_var; -- 
    end process;
    type_cast_4582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4582_inst_req_0;
      type_cast_4582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4582_inst_req_1;
      type_cast_4582_inst_ack_1<= rack(0);
      type_cast_4582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4581_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_4583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4586_inst
    process(conv66_4583) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv66_4583(31 downto 0);
      type_cast_4586_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4588_inst
    process(conv54_4450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv54_4450(31 downto 0);
      type_cast_4588_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4599_inst
    process(conv66_4583) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv66_4583(31 downto 0);
      type_cast_4599_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4601_inst
    process(add78_4499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add78_4499(31 downto 0);
      type_cast_4601_wire <= tmp_var; -- 
    end process;
    type_cast_4619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4619_inst_req_0;
      type_cast_4619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4619_inst_req_1;
      type_cast_4619_inst_ack_1<= rack(0);
      type_cast_4619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4618_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_4620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4624_inst_req_0;
      type_cast_4624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4624_inst_req_1;
      type_cast_4624_inst_ack_1<= rack(0);
      type_cast_4624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4623_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_4625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4648_inst
    process(add95_4645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add95_4645(31 downto 0);
      type_cast_4648_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4653_inst
    process(ASHR_i32_i32_4652_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4652_wire(31 downto 0);
      shr_4654 <= tmp_var; -- 
    end process;
    type_cast_4658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4658_inst_req_0;
      type_cast_4658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4658_inst_req_1;
      type_cast_4658_inst_ack_1<= rack(0);
      type_cast_4658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4657_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_4659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4677_inst_req_0;
      type_cast_4677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4677_inst_req_1;
      type_cast_4677_inst_ack_1<= rack(0);
      type_cast_4677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4676_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_4678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4731_inst
    process(add116_4708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add116_4708(31 downto 0);
      type_cast_4731_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4736_inst
    process(ASHR_i32_i32_4735_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4735_wire(31 downto 0);
      shr134_4737 <= tmp_var; -- 
    end process;
    type_cast_4741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4741_inst_req_0;
      type_cast_4741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4741_inst_req_1;
      type_cast_4741_inst_ack_1<= rack(0);
      type_cast_4741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4740_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom135_4742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4756_inst
    process(add132_4728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add132_4728(31 downto 0);
      type_cast_4756_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4761_inst
    process(ASHR_i32_i32_4760_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4760_wire(31 downto 0);
      shr139_4762 <= tmp_var; -- 
    end process;
    type_cast_4766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4766_inst_req_0;
      type_cast_4766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4766_inst_req_1;
      type_cast_4766_inst_ack_1<= rack(0);
      type_cast_4766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4765_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom140_4767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4784_inst_req_0;
      type_cast_4784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4784_inst_req_1;
      type_cast_4784_inst_ack_1<= rack(0);
      type_cast_4784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4783_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_4785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4794_inst
    process(add145_4791) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add145_4791(31 downto 0);
      type_cast_4794_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4796_inst
    process(conv36_4429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_4429(31 downto 0);
      type_cast_4796_wire <= tmp_var; -- 
    end process;
    type_cast_4823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4823_inst_req_0;
      type_cast_4823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4823_inst_req_1;
      type_cast_4823_inst_ack_1<= rack(0);
      type_cast_4823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4822_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_4824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4832_inst_req_0;
      type_cast_4832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4832_inst_req_1;
      type_cast_4832_inst_ack_1<= rack(0);
      type_cast_4832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp164_4829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc169_4833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4848_inst_req_0;
      type_cast_4848_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4848_inst_req_1;
      type_cast_4848_inst_ack_1<= rack(0);
      type_cast_4848_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4848_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4847_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv172_4849,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4868_inst_req_0;
      type_cast_4868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4868_inst_req_1;
      type_cast_4868_inst_ack_1<= rack(0);
      type_cast_4868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add153_4811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4868_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4872_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4872_inst_req_0;
      type_cast_4872_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4872_inst_req_1;
      type_cast_4872_inst_ack_1<= rack(0);
      type_cast_4872_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4872_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_4529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4872_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4874_inst_req_0;
      type_cast_4874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4874_inst_req_1;
      type_cast_4874_inst_ack_1<= rack(0);
      type_cast_4874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc169x_xix_x2_4838,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4874_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4878_inst_req_0;
      type_cast_4878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4878_inst_req_1;
      type_cast_4878_inst_ack_1<= rack(0);
      type_cast_4878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4878_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_4535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4878_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4880_inst_req_0;
      type_cast_4880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4880_inst_req_1;
      type_cast_4880_inst_ack_1<= rack(0);
      type_cast_4880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_4844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4880_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_4664_index_1_rename
    process(R_idxprom_4663_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_4663_resized;
      ov(13 downto 0) := iv;
      R_idxprom_4663_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4664_index_1_resize
    process(idxprom_4659) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_4659;
      ov := iv(13 downto 0);
      R_idxprom_4663_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4664_root_address_inst
    process(array_obj_ref_4664_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4664_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4664_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4747_index_1_rename
    process(R_idxprom135_4746_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom135_4746_resized;
      ov(13 downto 0) := iv;
      R_idxprom135_4746_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4747_index_1_resize
    process(idxprom135_4742) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom135_4742;
      ov := iv(13 downto 0);
      R_idxprom135_4746_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4747_root_address_inst
    process(array_obj_ref_4747_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4747_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4747_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4772_index_1_rename
    process(R_idxprom140_4771_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom140_4771_resized;
      ov(13 downto 0) := iv;
      R_idxprom140_4771_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4772_index_1_resize
    process(idxprom140_4767) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom140_4767;
      ov := iv(13 downto 0);
      R_idxprom140_4771_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4772_root_address_inst
    process(array_obj_ref_4772_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4772_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4772_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4668_addr_0
    process(ptr_deref_4668_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4668_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4668_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4668_base_resize
    process(arrayidx_4666) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_4666;
      ov := iv(13 downto 0);
      ptr_deref_4668_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4668_gather_scatter
    process(type_cast_4670_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_4670_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_4668_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4668_root_address_inst
    process(ptr_deref_4668_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4668_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4668_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4752_addr_0
    process(ptr_deref_4752_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4752_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4752_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4752_base_resize
    process(arrayidx136_4749) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx136_4749;
      ov := iv(13 downto 0);
      ptr_deref_4752_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4752_gather_scatter
    process(ptr_deref_4752_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4752_data_0;
      ov(63 downto 0) := iv;
      tmp137_4753 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4752_root_address_inst
    process(ptr_deref_4752_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4752_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4752_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4776_addr_0
    process(ptr_deref_4776_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4776_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4776_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4776_base_resize
    process(arrayidx141_4774) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx141_4774;
      ov := iv(13 downto 0);
      ptr_deref_4776_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4776_gather_scatter
    process(tmp137_4753) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp137_4753;
      ov(63 downto 0) := iv;
      ptr_deref_4776_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4776_root_address_inst
    process(ptr_deref_4776_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4776_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4776_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_4572_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_4571;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4572_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4572_branch_req_0,
          ack0 => if_stmt_4572_branch_ack_0,
          ack1 => if_stmt_4572_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4609_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond193_4608;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4609_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4609_branch_req_0,
          ack0 => if_stmt_4609_branch_ack_0,
          ack1 => if_stmt_4609_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4799_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp148_4798;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4799_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4799_branch_req_0,
          ack0 => if_stmt_4799_branch_ack_0,
          ack1 => if_stmt_4799_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4855_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp179_4854;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4855_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4855_branch_req_0,
          ack0 => if_stmt_4855_branch_ack_0,
          ack1 => if_stmt_4855_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_4810_inst
    process(kx_x1_4522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_4522, type_cast_4809_wire_constant, tmp_var);
      add153_4811 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4818_inst
    process(jx_x1_4535) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_4535, type_cast_4817_wire_constant, tmp_var);
      inc_4819 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4837_inst
    process(inc169_4833, ix_x2_4529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc169_4833, ix_x2_4529, tmp_var);
      inc169x_xix_x2_4838 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4479_inst
    process(shl_4475, conv38_4433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_4475, conv38_4433, tmp_var);
      add163_4480 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4488_inst
    process(shl_4475, conv174_4484) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_4475, conv174_4484, tmp_var);
      add178_4489 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4493_inst
    process(conv54_4450, conv174_4484) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv54_4450, conv174_4484, tmp_var);
      add_4494 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4498_inst
    process(conv54_4450, conv38_4433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv54_4450, conv38_4433, tmp_var);
      add78_4499 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4639_inst
    process(mul94_4635, conv83_4620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul94_4635, conv83_4620, tmp_var);
      add89_4640 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4644_inst
    process(add89_4640, mul88_4630) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add89_4640, mul88_4630, tmp_var);
      add95_4645 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4702_inst
    process(mul115_4698, conv99_4678) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul115_4698, conv99_4678, tmp_var);
      add107_4703 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4707_inst
    process(add107_4703, mul106_4688) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add107_4703, mul106_4688, tmp_var);
      add116_4708 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4722_inst
    process(mul131_4718, conv99_4678) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul131_4718, conv99_4678, tmp_var);
      add126_4723 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4727_inst
    process(add126_4723, mul125_4713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add126_4723, mul125_4713, tmp_var);
      add132_4728 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4790_inst
    process(conv144_4785) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv144_4785, type_cast_4789_wire_constant, tmp_var);
      add145_4791 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_4570_inst
    process(cmpx_xnot_4559, cmp62_4566) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_4559, cmp62_4566, tmp_var);
      orx_xcond_4571 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_4607_inst
    process(cmp69x_xnot_4596, cmp79_4603) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp69x_xnot_4596, cmp79_4603, tmp_var);
      orx_xcond193_4608 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4467_inst
    process(type_cast_4463_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4463_wire, type_cast_4466_wire_constant, tmp_var);
      ASHR_i32_i32_4467_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4517_inst
    process(type_cast_4513_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4513_wire, type_cast_4516_wire_constant, tmp_var);
      ASHR_i32_i32_4517_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4652_inst
    process(type_cast_4648_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4648_wire, type_cast_4651_wire_constant, tmp_var);
      ASHR_i32_i32_4652_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4735_inst
    process(type_cast_4731_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4731_wire, type_cast_4734_wire_constant, tmp_var);
      ASHR_i32_i32_4735_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4760_inst
    process(type_cast_4756_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4756_wire, type_cast_4759_wire_constant, tmp_var);
      ASHR_i32_i32_4760_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4828_inst
    process(conv158_4824, add163_4480) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv158_4824, add163_4480, tmp_var);
      cmp164_4829 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4853_inst
    process(conv172_4849, add178_4489) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv172_4849, add178_4489, tmp_var);
      cmp179_4854 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4408_inst
    process(conv_4403) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_4403, type_cast_4407_wire_constant, tmp_var);
      div_4409 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4424_inst
    process(mul_4419) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul_4419, type_cast_4423_wire_constant, tmp_var);
      div11_4425 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_4418_inst
    process(conv10_4413) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv10_4413, type_cast_4417_wire_constant, tmp_var);
      mul_4419 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4445_inst
    process(conv43_4437, conv45_4441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv43_4437, conv45_4441, tmp_var);
      mul46_4446 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4509_inst
    process(mul39_4505, conv36_4429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul39_4505, conv36_4429, tmp_var);
      sext_4510 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4629_inst
    process(conv87_4625, conv85_4454) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv87_4625, conv85_4454, tmp_var);
      mul88_4630 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4634_inst
    process(conv52_4546, conv91_4469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv52_4546, conv91_4469, tmp_var);
      mul94_4635 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4687_inst
    process(sub_4683, conv36_4429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_4683, conv36_4429, tmp_var);
      mul106_4688 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4697_inst
    process(sub114_4693, conv109_4519) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub114_4693, conv109_4519, tmp_var);
      mul115_4698 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4712_inst
    process(conv66_4583, conv85_4454) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv66_4583, conv85_4454, tmp_var);
      mul125_4713 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4717_inst
    process(conv52_4546, conv91_4469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv52_4546, conv91_4469, tmp_var);
      mul131_4718 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4459_inst
    process(mul46_4446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul46_4446, type_cast_4458_wire_constant, tmp_var);
      sext192_4460 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4474_inst
    process(conv54_4450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv54_4450, type_cast_4473_wire_constant, tmp_var);
      shl_4475 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4504_inst
    process(conv38_4433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv38_4433, type_cast_4503_wire_constant, tmp_var);
      mul39_4505 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4552_inst
    process(type_cast_4549_wire, type_cast_4551_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4549_wire, type_cast_4551_wire, tmp_var);
      cmp_4553 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4565_inst
    process(type_cast_4562_wire, type_cast_4564_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4562_wire, type_cast_4564_wire, tmp_var);
      cmp62_4566 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4589_inst
    process(type_cast_4586_wire, type_cast_4588_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4586_wire, type_cast_4588_wire, tmp_var);
      cmp69_4590 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4602_inst
    process(type_cast_4599_wire, type_cast_4601_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4599_wire, type_cast_4601_wire, tmp_var);
      cmp79_4603 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4797_inst
    process(type_cast_4794_wire, type_cast_4796_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4794_wire, type_cast_4796_wire, tmp_var);
      cmp148_4798 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4682_inst
    process(conv66_4583, conv54_4450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv66_4583, conv54_4450, tmp_var);
      sub_4683 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4692_inst
    process(conv52_4546, conv54_4450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv52_4546, conv54_4450, tmp_var);
      sub114_4693 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_4558_inst
    process(cmp_4553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_4553, type_cast_4557_wire_constant, tmp_var);
      cmpx_xnot_4559 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_4595_inst
    process(cmp69_4590) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp69_4590, type_cast_4594_wire_constant, tmp_var);
      cmp69x_xnot_4596 <= tmp_var; --
    end process;
    -- shared split operator group (46) : array_obj_ref_4664_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_4663_scaled;
      array_obj_ref_4664_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4664_index_offset_req_0;
      array_obj_ref_4664_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4664_index_offset_req_1;
      array_obj_ref_4664_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_4747_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom135_4746_scaled;
      array_obj_ref_4747_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4747_index_offset_req_0;
      array_obj_ref_4747_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4747_index_offset_req_1;
      array_obj_ref_4747_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_4772_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom140_4771_scaled;
      array_obj_ref_4772_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4772_index_offset_req_0;
      array_obj_ref_4772_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4772_index_offset_req_1;
      array_obj_ref_4772_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- unary operator type_cast_4544_inst
    process(ix_x2_4529) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_4529, tmp_var);
      type_cast_4544_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4581_inst
    process(jx_x1_4535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_4535, tmp_var);
      type_cast_4581_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4618_inst
    process(kx_x1_4522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_4522, tmp_var);
      type_cast_4618_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4623_inst
    process(jx_x1_4535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_4535, tmp_var);
      type_cast_4623_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4657_inst
    process(shr_4654) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_4654, tmp_var);
      type_cast_4657_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4676_inst
    process(kx_x1_4522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_4522, tmp_var);
      type_cast_4676_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4740_inst
    process(shr134_4737) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr134_4737, tmp_var);
      type_cast_4740_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4765_inst
    process(shr139_4762) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr139_4762, tmp_var);
      type_cast_4765_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4783_inst
    process(kx_x1_4522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_4522, tmp_var);
      type_cast_4783_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4822_inst
    process(inc_4819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_4819, tmp_var);
      type_cast_4822_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4847_inst
    process(inc169x_xix_x2_4838) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc169x_xix_x2_4838, tmp_var);
      type_cast_4847_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_4752_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_4752_load_0_req_0;
      ptr_deref_4752_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_4752_load_0_req_1;
      ptr_deref_4752_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_4752_word_address_0;
      ptr_deref_4752_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_4776_store_0 ptr_deref_4668_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_4776_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4668_store_0_req_0;
      ptr_deref_4776_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4668_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_4776_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4668_store_0_req_1;
      ptr_deref_4776_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4668_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_4776_word_address_0 & ptr_deref_4668_word_address_0;
      data_in <= ptr_deref_4776_data_0 & ptr_deref_4668_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 19,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block7_starting_4379_inst RPIPE_Block7_starting_4382_inst RPIPE_Block7_starting_4385_inst RPIPE_Block7_starting_4388_inst RPIPE_Block7_starting_4391_inst RPIPE_Block7_starting_4394_inst RPIPE_Block7_starting_4397_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block7_starting_4379_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block7_starting_4382_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block7_starting_4385_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block7_starting_4388_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block7_starting_4391_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block7_starting_4394_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block7_starting_4397_inst_req_0;
      RPIPE_Block7_starting_4379_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block7_starting_4382_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block7_starting_4385_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block7_starting_4388_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block7_starting_4391_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block7_starting_4394_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block7_starting_4397_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block7_starting_4379_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block7_starting_4382_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block7_starting_4385_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block7_starting_4388_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block7_starting_4391_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block7_starting_4394_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block7_starting_4397_inst_req_1;
      RPIPE_Block7_starting_4379_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block7_starting_4382_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block7_starting_4385_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block7_starting_4388_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block7_starting_4391_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block7_starting_4394_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block7_starting_4397_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call_4380 <= data_out(55 downto 48);
      call1_4383 <= data_out(47 downto 40);
      call2_4386 <= data_out(39 downto 32);
      call3_4389 <= data_out(31 downto 24);
      call4_4392 <= data_out(23 downto 16);
      call5_4395 <= data_out(15 downto 8);
      call6_4398 <= data_out(7 downto 0);
      Block7_starting_read_0_gI: SplitGuardInterface generic map(name => "Block7_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block7_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block7_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block7_starting_pipe_read_req(0),
          oack => Block7_starting_pipe_read_ack(0),
          odata => Block7_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block7_complete_4885_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block7_complete_4885_inst_req_0;
      WPIPE_Block7_complete_4885_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block7_complete_4885_inst_req_1;
      WPIPE_Block7_complete_4885_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_4887_wire_constant;
      Block7_complete_write_0_gI: SplitGuardInterface generic map(name => "Block7_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block7_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block7_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block7_complete_pipe_write_req(0),
          oack => Block7_complete_pipe_write_ack(0),
          odata => Block7_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_H_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(7 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(7 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(111 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(511 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(167 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(7 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(15 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(7 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(7 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(111 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(159 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(7 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(511 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_size :  std_logic_vector(31 downto 0);
  signal sendOutput_in_args    : std_logic_vector(31 downto 0);
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_data: std_logic_vector(31 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block3_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block4_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block4_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block4_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block5_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block5_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block5_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block6_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block6_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block6_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block7_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block7_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block7_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block3_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block7_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block7_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block7_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      Block4_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block4_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block4_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block5_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block5_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block5_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block6_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block6_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block6_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_data : out  std_logic_vector(31 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- declarations related to module zeropad3D_A
  component zeropad3D_A is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_A
  signal zeropad3D_A_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_A_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_A_start_req : std_logic;
  signal zeropad3D_A_start_ack : std_logic;
  signal zeropad3D_A_fin_req   : std_logic;
  signal zeropad3D_A_fin_ack : std_logic;
  -- declarations related to module zeropad3D_B
  component zeropad3D_B is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block1_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_B
  signal zeropad3D_B_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_B_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_B_start_req : std_logic;
  signal zeropad3D_B_start_ack : std_logic;
  signal zeropad3D_B_fin_req   : std_logic;
  signal zeropad3D_B_fin_ack : std_logic;
  -- declarations related to module zeropad3D_C
  component zeropad3D_C is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block2_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_C
  signal zeropad3D_C_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_C_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_C_start_req : std_logic;
  signal zeropad3D_C_start_ack : std_logic;
  signal zeropad3D_C_fin_req   : std_logic;
  signal zeropad3D_C_fin_ack : std_logic;
  -- declarations related to module zeropad3D_D
  component zeropad3D_D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block3_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block3_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_D
  signal zeropad3D_D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_D_start_req : std_logic;
  signal zeropad3D_D_start_ack : std_logic;
  signal zeropad3D_D_fin_req   : std_logic;
  signal zeropad3D_D_fin_ack : std_logic;
  -- declarations related to module zeropad3D_E
  component zeropad3D_E is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block4_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block4_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block4_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block4_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block4_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block4_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_E
  signal zeropad3D_E_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_E_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_E_start_req : std_logic;
  signal zeropad3D_E_start_ack : std_logic;
  signal zeropad3D_E_fin_req   : std_logic;
  signal zeropad3D_E_fin_ack : std_logic;
  -- declarations related to module zeropad3D_F
  component zeropad3D_F is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block5_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block5_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block5_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block5_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block5_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block5_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_F
  signal zeropad3D_F_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_F_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_F_start_req : std_logic;
  signal zeropad3D_F_start_ack : std_logic;
  signal zeropad3D_F_fin_req   : std_logic;
  signal zeropad3D_F_fin_ack : std_logic;
  -- declarations related to module zeropad3D_G
  component zeropad3D_G is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block6_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block6_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block6_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block6_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block6_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block6_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_G
  signal zeropad3D_G_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_G_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_G_start_req : std_logic;
  signal zeropad3D_G_start_ack : std_logic;
  signal zeropad3D_G_fin_req   : std_logic;
  signal zeropad3D_G_fin_ack : std_logic;
  -- declarations related to module zeropad3D_H
  component zeropad3D_H is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block7_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block7_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block7_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block7_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block7_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block7_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_H
  signal zeropad3D_H_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_H_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_H_start_req : std_logic;
  signal zeropad3D_H_start_ack : std_logic;
  signal zeropad3D_H_fin_req   : std_logic;
  signal zeropad3D_H_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_complete
  signal Block0_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_complete
  signal Block0_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_starting
  signal Block0_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_starting
  signal Block0_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_complete
  signal Block1_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block1_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_complete
  signal Block1_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block1_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_starting
  signal Block1_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block1_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_starting
  signal Block1_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block1_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_complete
  signal Block2_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block2_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_complete
  signal Block2_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block2_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_starting
  signal Block2_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block2_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_starting
  signal Block2_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block2_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_complete
  signal Block3_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block3_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_complete
  signal Block3_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block3_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_starting
  signal Block3_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block3_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_starting
  signal Block3_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block3_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block4_complete
  signal Block4_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block4_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block4_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block4_complete
  signal Block4_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block4_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block4_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block4_starting
  signal Block4_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block4_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block4_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block4_starting
  signal Block4_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block4_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block4_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block5_complete
  signal Block5_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block5_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block5_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block5_complete
  signal Block5_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block5_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block5_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block5_starting
  signal Block5_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block5_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block5_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block5_starting
  signal Block5_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block5_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block5_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block6_complete
  signal Block6_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block6_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block6_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block6_complete
  signal Block6_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block6_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block6_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block6_starting
  signal Block6_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block6_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block6_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block6_starting
  signal Block6_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block6_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block6_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block7_complete
  signal Block7_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block7_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block7_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block7_complete
  signal Block7_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block7_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block7_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block7_starting
  signal Block7_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block7_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block7_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block7_starting
  signal Block7_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block7_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block7_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  sendOutput_size <= sendOutput_in_args(31 downto 0);
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_data  => sendOutput_call_data,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      call_mdata => sendOutput_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendOutput_size,
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(20 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(0 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      Block0_complete_pipe_read_req => Block0_complete_pipe_read_req(0 downto 0),
      Block0_complete_pipe_read_ack => Block0_complete_pipe_read_ack(0 downto 0),
      Block0_complete_pipe_read_data => Block0_complete_pipe_read_data(7 downto 0),
      Block1_complete_pipe_read_req => Block1_complete_pipe_read_req(0 downto 0),
      Block1_complete_pipe_read_ack => Block1_complete_pipe_read_ack(0 downto 0),
      Block1_complete_pipe_read_data => Block1_complete_pipe_read_data(7 downto 0),
      Block3_complete_pipe_read_req => Block3_complete_pipe_read_req(0 downto 0),
      Block3_complete_pipe_read_ack => Block3_complete_pipe_read_ack(0 downto 0),
      Block3_complete_pipe_read_data => Block3_complete_pipe_read_data(7 downto 0),
      Block4_complete_pipe_read_req => Block4_complete_pipe_read_req(0 downto 0),
      Block4_complete_pipe_read_ack => Block4_complete_pipe_read_ack(0 downto 0),
      Block4_complete_pipe_read_data => Block4_complete_pipe_read_data(7 downto 0),
      Block2_complete_pipe_read_req => Block2_complete_pipe_read_req(0 downto 0),
      Block2_complete_pipe_read_ack => Block2_complete_pipe_read_ack(0 downto 0),
      Block2_complete_pipe_read_data => Block2_complete_pipe_read_data(7 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      Block5_complete_pipe_read_req => Block5_complete_pipe_read_req(0 downto 0),
      Block5_complete_pipe_read_ack => Block5_complete_pipe_read_ack(0 downto 0),
      Block5_complete_pipe_read_data => Block5_complete_pipe_read_data(7 downto 0),
      Block6_complete_pipe_read_req => Block6_complete_pipe_read_req(0 downto 0),
      Block6_complete_pipe_read_ack => Block6_complete_pipe_read_ack(0 downto 0),
      Block6_complete_pipe_read_data => Block6_complete_pipe_read_data(7 downto 0),
      Block7_complete_pipe_read_req => Block7_complete_pipe_read_req(0 downto 0),
      Block7_complete_pipe_read_ack => Block7_complete_pipe_read_ack(0 downto 0),
      Block7_complete_pipe_read_data => Block7_complete_pipe_read_data(7 downto 0),
      Block1_starting_pipe_write_req => Block1_starting_pipe_write_req(0 downto 0),
      Block1_starting_pipe_write_ack => Block1_starting_pipe_write_ack(0 downto 0),
      Block1_starting_pipe_write_data => Block1_starting_pipe_write_data(7 downto 0),
      Block0_starting_pipe_write_req => Block0_starting_pipe_write_req(0 downto 0),
      Block0_starting_pipe_write_ack => Block0_starting_pipe_write_ack(0 downto 0),
      Block0_starting_pipe_write_data => Block0_starting_pipe_write_data(7 downto 0),
      Block3_starting_pipe_write_req => Block3_starting_pipe_write_req(0 downto 0),
      Block3_starting_pipe_write_ack => Block3_starting_pipe_write_ack(0 downto 0),
      Block3_starting_pipe_write_data => Block3_starting_pipe_write_data(7 downto 0),
      Block2_starting_pipe_write_req => Block2_starting_pipe_write_req(0 downto 0),
      Block2_starting_pipe_write_ack => Block2_starting_pipe_write_ack(0 downto 0),
      Block2_starting_pipe_write_data => Block2_starting_pipe_write_data(7 downto 0),
      Block7_starting_pipe_write_req => Block7_starting_pipe_write_req(0 downto 0),
      Block7_starting_pipe_write_ack => Block7_starting_pipe_write_ack(0 downto 0),
      Block7_starting_pipe_write_data => Block7_starting_pipe_write_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      Block4_starting_pipe_write_req => Block4_starting_pipe_write_req(0 downto 0),
      Block4_starting_pipe_write_ack => Block4_starting_pipe_write_ack(0 downto 0),
      Block4_starting_pipe_write_data => Block4_starting_pipe_write_data(7 downto 0),
      Block5_starting_pipe_write_req => Block5_starting_pipe_write_req(0 downto 0),
      Block5_starting_pipe_write_ack => Block5_starting_pipe_write_ack(0 downto 0),
      Block5_starting_pipe_write_data => Block5_starting_pipe_write_data(7 downto 0),
      Block6_starting_pipe_write_req => Block6_starting_pipe_write_req(0 downto 0),
      Block6_starting_pipe_write_ack => Block6_starting_pipe_write_ack(0 downto 0),
      Block6_starting_pipe_write_data => Block6_starting_pipe_write_data(7 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_data => sendOutput_call_data(31 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  -- module zeropad3D_A
  zeropad3D_A_instance:zeropad3D_A-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_A_start_req,
      start_ack => zeropad3D_A_start_ack,
      fin_req => zeropad3D_A_fin_req,
      fin_ack => zeropad3D_A_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(7 downto 7),
      memory_space_1_lr_ack => memory_space_1_lr_ack(7 downto 7),
      memory_space_1_lr_addr => memory_space_1_lr_addr(111 downto 98),
      memory_space_1_lr_tag => memory_space_1_lr_tag(159 downto 140),
      memory_space_1_lc_req => memory_space_1_lc_req(7 downto 7),
      memory_space_1_lc_ack => memory_space_1_lc_ack(7 downto 7),
      memory_space_1_lc_data => memory_space_1_lc_data(511 downto 448),
      memory_space_1_lc_tag => memory_space_1_lc_tag(7 downto 7),
      memory_space_0_sr_req => memory_space_0_sr_req(7 downto 7),
      memory_space_0_sr_ack => memory_space_0_sr_ack(7 downto 7),
      memory_space_0_sr_addr => memory_space_0_sr_addr(111 downto 98),
      memory_space_0_sr_data => memory_space_0_sr_data(511 downto 448),
      memory_space_0_sr_tag => memory_space_0_sr_tag(167 downto 147),
      memory_space_0_sc_req => memory_space_0_sc_req(7 downto 7),
      memory_space_0_sc_ack => memory_space_0_sc_ack(7 downto 7),
      memory_space_0_sc_tag => memory_space_0_sc_tag(15 downto 14),
      Block0_starting_pipe_read_req => Block0_starting_pipe_read_req(0 downto 0),
      Block0_starting_pipe_read_ack => Block0_starting_pipe_read_ack(0 downto 0),
      Block0_starting_pipe_read_data => Block0_starting_pipe_read_data(7 downto 0),
      Block0_complete_pipe_write_req => Block0_complete_pipe_write_req(0 downto 0),
      Block0_complete_pipe_write_ack => Block0_complete_pipe_write_ack(0 downto 0),
      Block0_complete_pipe_write_data => Block0_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_A_tag_in,
      tag_out => zeropad3D_A_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_A_tag_in <= (others => '0');
  zeropad3D_A_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_A_start_req, start_ack => zeropad3D_A_start_ack,  fin_req => zeropad3D_A_fin_req,  fin_ack => zeropad3D_A_fin_ack);
  -- module zeropad3D_B
  zeropad3D_B_instance:zeropad3D_B-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_B_start_req,
      start_ack => zeropad3D_B_start_ack,
      fin_req => zeropad3D_B_fin_req,
      fin_ack => zeropad3D_B_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(6 downto 6),
      memory_space_1_lr_ack => memory_space_1_lr_ack(6 downto 6),
      memory_space_1_lr_addr => memory_space_1_lr_addr(97 downto 84),
      memory_space_1_lr_tag => memory_space_1_lr_tag(139 downto 120),
      memory_space_1_lc_req => memory_space_1_lc_req(6 downto 6),
      memory_space_1_lc_ack => memory_space_1_lc_ack(6 downto 6),
      memory_space_1_lc_data => memory_space_1_lc_data(447 downto 384),
      memory_space_1_lc_tag => memory_space_1_lc_tag(6 downto 6),
      memory_space_0_sr_req => memory_space_0_sr_req(6 downto 6),
      memory_space_0_sr_ack => memory_space_0_sr_ack(6 downto 6),
      memory_space_0_sr_addr => memory_space_0_sr_addr(97 downto 84),
      memory_space_0_sr_data => memory_space_0_sr_data(447 downto 384),
      memory_space_0_sr_tag => memory_space_0_sr_tag(146 downto 126),
      memory_space_0_sc_req => memory_space_0_sc_req(6 downto 6),
      memory_space_0_sc_ack => memory_space_0_sc_ack(6 downto 6),
      memory_space_0_sc_tag => memory_space_0_sc_tag(13 downto 12),
      Block1_starting_pipe_read_req => Block1_starting_pipe_read_req(0 downto 0),
      Block1_starting_pipe_read_ack => Block1_starting_pipe_read_ack(0 downto 0),
      Block1_starting_pipe_read_data => Block1_starting_pipe_read_data(7 downto 0),
      Block1_complete_pipe_write_req => Block1_complete_pipe_write_req(0 downto 0),
      Block1_complete_pipe_write_ack => Block1_complete_pipe_write_ack(0 downto 0),
      Block1_complete_pipe_write_data => Block1_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_B_tag_in,
      tag_out => zeropad3D_B_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_B_tag_in <= (others => '0');
  zeropad3D_B_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_B_start_req, start_ack => zeropad3D_B_start_ack,  fin_req => zeropad3D_B_fin_req,  fin_ack => zeropad3D_B_fin_ack);
  -- module zeropad3D_C
  zeropad3D_C_instance:zeropad3D_C-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_C_start_req,
      start_ack => zeropad3D_C_start_ack,
      fin_req => zeropad3D_C_fin_req,
      fin_ack => zeropad3D_C_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(5 downto 5),
      memory_space_1_lr_ack => memory_space_1_lr_ack(5 downto 5),
      memory_space_1_lr_addr => memory_space_1_lr_addr(83 downto 70),
      memory_space_1_lr_tag => memory_space_1_lr_tag(119 downto 100),
      memory_space_1_lc_req => memory_space_1_lc_req(5 downto 5),
      memory_space_1_lc_ack => memory_space_1_lc_ack(5 downto 5),
      memory_space_1_lc_data => memory_space_1_lc_data(383 downto 320),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 5),
      memory_space_0_sr_req => memory_space_0_sr_req(5 downto 5),
      memory_space_0_sr_ack => memory_space_0_sr_ack(5 downto 5),
      memory_space_0_sr_addr => memory_space_0_sr_addr(83 downto 70),
      memory_space_0_sr_data => memory_space_0_sr_data(383 downto 320),
      memory_space_0_sr_tag => memory_space_0_sr_tag(125 downto 105),
      memory_space_0_sc_req => memory_space_0_sc_req(5 downto 5),
      memory_space_0_sc_ack => memory_space_0_sc_ack(5 downto 5),
      memory_space_0_sc_tag => memory_space_0_sc_tag(11 downto 10),
      Block2_starting_pipe_read_req => Block2_starting_pipe_read_req(0 downto 0),
      Block2_starting_pipe_read_ack => Block2_starting_pipe_read_ack(0 downto 0),
      Block2_starting_pipe_read_data => Block2_starting_pipe_read_data(7 downto 0),
      Block2_complete_pipe_write_req => Block2_complete_pipe_write_req(0 downto 0),
      Block2_complete_pipe_write_ack => Block2_complete_pipe_write_ack(0 downto 0),
      Block2_complete_pipe_write_data => Block2_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_C_tag_in,
      tag_out => zeropad3D_C_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_C_tag_in <= (others => '0');
  zeropad3D_C_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_C_start_req, start_ack => zeropad3D_C_start_ack,  fin_req => zeropad3D_C_fin_req,  fin_ack => zeropad3D_C_fin_ack);
  -- module zeropad3D_D
  zeropad3D_D_instance:zeropad3D_D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_D_start_req,
      start_ack => zeropad3D_D_start_ack,
      fin_req => zeropad3D_D_fin_req,
      fin_ack => zeropad3D_D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(69 downto 56),
      memory_space_1_lr_tag => memory_space_1_lr_tag(99 downto 80),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(319 downto 256),
      memory_space_1_lc_tag => memory_space_1_lc_tag(4 downto 4),
      memory_space_0_sr_req => memory_space_0_sr_req(4 downto 4),
      memory_space_0_sr_ack => memory_space_0_sr_ack(4 downto 4),
      memory_space_0_sr_addr => memory_space_0_sr_addr(69 downto 56),
      memory_space_0_sr_data => memory_space_0_sr_data(319 downto 256),
      memory_space_0_sr_tag => memory_space_0_sr_tag(104 downto 84),
      memory_space_0_sc_req => memory_space_0_sc_req(4 downto 4),
      memory_space_0_sc_ack => memory_space_0_sc_ack(4 downto 4),
      memory_space_0_sc_tag => memory_space_0_sc_tag(9 downto 8),
      Block3_starting_pipe_read_req => Block3_starting_pipe_read_req(0 downto 0),
      Block3_starting_pipe_read_ack => Block3_starting_pipe_read_ack(0 downto 0),
      Block3_starting_pipe_read_data => Block3_starting_pipe_read_data(7 downto 0),
      Block3_complete_pipe_write_req => Block3_complete_pipe_write_req(0 downto 0),
      Block3_complete_pipe_write_ack => Block3_complete_pipe_write_ack(0 downto 0),
      Block3_complete_pipe_write_data => Block3_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_D_tag_in,
      tag_out => zeropad3D_D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_D_tag_in <= (others => '0');
  zeropad3D_D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_D_start_req, start_ack => zeropad3D_D_start_ack,  fin_req => zeropad3D_D_fin_req,  fin_ack => zeropad3D_D_fin_ack);
  -- module zeropad3D_E
  zeropad3D_E_instance:zeropad3D_E-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_E_start_req,
      start_ack => zeropad3D_E_start_ack,
      fin_req => zeropad3D_E_fin_req,
      fin_ack => zeropad3D_E_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(79 downto 60),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_0_sr_req => memory_space_0_sr_req(3 downto 3),
      memory_space_0_sr_ack => memory_space_0_sr_ack(3 downto 3),
      memory_space_0_sr_addr => memory_space_0_sr_addr(55 downto 42),
      memory_space_0_sr_data => memory_space_0_sr_data(255 downto 192),
      memory_space_0_sr_tag => memory_space_0_sr_tag(83 downto 63),
      memory_space_0_sc_req => memory_space_0_sc_req(3 downto 3),
      memory_space_0_sc_ack => memory_space_0_sc_ack(3 downto 3),
      memory_space_0_sc_tag => memory_space_0_sc_tag(7 downto 6),
      Block4_starting_pipe_read_req => Block4_starting_pipe_read_req(0 downto 0),
      Block4_starting_pipe_read_ack => Block4_starting_pipe_read_ack(0 downto 0),
      Block4_starting_pipe_read_data => Block4_starting_pipe_read_data(7 downto 0),
      Block4_complete_pipe_write_req => Block4_complete_pipe_write_req(0 downto 0),
      Block4_complete_pipe_write_ack => Block4_complete_pipe_write_ack(0 downto 0),
      Block4_complete_pipe_write_data => Block4_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_E_tag_in,
      tag_out => zeropad3D_E_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_E_tag_in <= (others => '0');
  zeropad3D_E_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_E_start_req, start_ack => zeropad3D_E_start_ack,  fin_req => zeropad3D_E_fin_req,  fin_ack => zeropad3D_E_fin_ack);
  -- module zeropad3D_F
  zeropad3D_F_instance:zeropad3D_F-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_F_start_req,
      start_ack => zeropad3D_F_start_ack,
      fin_req => zeropad3D_F_fin_req,
      fin_ack => zeropad3D_F_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(59 downto 40),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_0_sr_req => memory_space_0_sr_req(2 downto 2),
      memory_space_0_sr_ack => memory_space_0_sr_ack(2 downto 2),
      memory_space_0_sr_addr => memory_space_0_sr_addr(41 downto 28),
      memory_space_0_sr_data => memory_space_0_sr_data(191 downto 128),
      memory_space_0_sr_tag => memory_space_0_sr_tag(62 downto 42),
      memory_space_0_sc_req => memory_space_0_sc_req(2 downto 2),
      memory_space_0_sc_ack => memory_space_0_sc_ack(2 downto 2),
      memory_space_0_sc_tag => memory_space_0_sc_tag(5 downto 4),
      Block5_starting_pipe_read_req => Block5_starting_pipe_read_req(0 downto 0),
      Block5_starting_pipe_read_ack => Block5_starting_pipe_read_ack(0 downto 0),
      Block5_starting_pipe_read_data => Block5_starting_pipe_read_data(7 downto 0),
      Block5_complete_pipe_write_req => Block5_complete_pipe_write_req(0 downto 0),
      Block5_complete_pipe_write_ack => Block5_complete_pipe_write_ack(0 downto 0),
      Block5_complete_pipe_write_data => Block5_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_F_tag_in,
      tag_out => zeropad3D_F_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_F_tag_in <= (others => '0');
  zeropad3D_F_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_F_start_req, start_ack => zeropad3D_F_start_ack,  fin_req => zeropad3D_F_fin_req,  fin_ack => zeropad3D_F_fin_ack);
  -- module zeropad3D_G
  zeropad3D_G_instance:zeropad3D_G-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_G_start_req,
      start_ack => zeropad3D_G_start_ack,
      fin_req => zeropad3D_G_fin_req,
      fin_ack => zeropad3D_G_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(39 downto 20),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(27 downto 14),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(41 downto 21),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      Block6_starting_pipe_read_req => Block6_starting_pipe_read_req(0 downto 0),
      Block6_starting_pipe_read_ack => Block6_starting_pipe_read_ack(0 downto 0),
      Block6_starting_pipe_read_data => Block6_starting_pipe_read_data(7 downto 0),
      Block6_complete_pipe_write_req => Block6_complete_pipe_write_req(0 downto 0),
      Block6_complete_pipe_write_ack => Block6_complete_pipe_write_ack(0 downto 0),
      Block6_complete_pipe_write_data => Block6_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_G_tag_in,
      tag_out => zeropad3D_G_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_G_tag_in <= (others => '0');
  zeropad3D_G_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_G_start_req, start_ack => zeropad3D_G_start_ack,  fin_req => zeropad3D_G_fin_req,  fin_ack => zeropad3D_G_fin_ack);
  -- module zeropad3D_H
  zeropad3D_H_instance:zeropad3D_H-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_H_start_req,
      start_ack => zeropad3D_H_start_ack,
      fin_req => zeropad3D_H_fin_req,
      fin_ack => zeropad3D_H_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(20 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Block7_starting_pipe_read_req => Block7_starting_pipe_read_req(0 downto 0),
      Block7_starting_pipe_read_ack => Block7_starting_pipe_read_ack(0 downto 0),
      Block7_starting_pipe_read_data => Block7_starting_pipe_read_data(7 downto 0),
      Block7_complete_pipe_write_req => Block7_complete_pipe_write_req(0 downto 0),
      Block7_complete_pipe_write_ack => Block7_complete_pipe_write_ack(0 downto 0),
      Block7_complete_pipe_write_data => Block7_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_H_tag_in,
      tag_out => zeropad3D_H_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_H_tag_in <= (others => '0');
  zeropad3D_H_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_H_start_req, start_ack => zeropad3D_H_start_ack,  fin_req => zeropad3D_H_fin_req,  fin_ack => zeropad3D_H_fin_ack);
  Block0_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_complete_pipe_read_req,
      read_ack => Block0_complete_pipe_read_ack,
      read_data => Block0_complete_pipe_read_data,
      write_req => Block0_complete_pipe_write_req,
      write_ack => Block0_complete_pipe_write_ack,
      write_data => Block0_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_starting_pipe_read_req,
      read_ack => Block0_starting_pipe_read_ack,
      read_data => Block0_starting_pipe_read_data,
      write_req => Block0_starting_pipe_write_req,
      write_ack => Block0_starting_pipe_write_ack,
      write_data => Block0_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_complete_pipe_read_req,
      read_ack => Block1_complete_pipe_read_ack,
      read_data => Block1_complete_pipe_read_data,
      write_req => Block1_complete_pipe_write_req,
      write_ack => Block1_complete_pipe_write_ack,
      write_data => Block1_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_starting_pipe_read_req,
      read_ack => Block1_starting_pipe_read_ack,
      read_data => Block1_starting_pipe_read_data,
      write_req => Block1_starting_pipe_write_req,
      write_ack => Block1_starting_pipe_write_ack,
      write_data => Block1_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_complete_pipe_read_req,
      read_ack => Block2_complete_pipe_read_ack,
      read_data => Block2_complete_pipe_read_data,
      write_req => Block2_complete_pipe_write_req,
      write_ack => Block2_complete_pipe_write_ack,
      write_data => Block2_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_starting_pipe_read_req,
      read_ack => Block2_starting_pipe_read_ack,
      read_data => Block2_starting_pipe_read_data,
      write_req => Block2_starting_pipe_write_req,
      write_ack => Block2_starting_pipe_write_ack,
      write_data => Block2_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_complete_pipe_read_req,
      read_ack => Block3_complete_pipe_read_ack,
      read_data => Block3_complete_pipe_read_data,
      write_req => Block3_complete_pipe_write_req,
      write_ack => Block3_complete_pipe_write_ack,
      write_data => Block3_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_starting_pipe_read_req,
      read_ack => Block3_starting_pipe_read_ack,
      read_data => Block3_starting_pipe_read_data,
      write_req => Block3_starting_pipe_write_req,
      write_ack => Block3_starting_pipe_write_ack,
      write_data => Block3_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block4_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block4_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block4_complete_pipe_read_req,
      read_ack => Block4_complete_pipe_read_ack,
      read_data => Block4_complete_pipe_read_data,
      write_req => Block4_complete_pipe_write_req,
      write_ack => Block4_complete_pipe_write_ack,
      write_data => Block4_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block4_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block4_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block4_starting_pipe_read_req,
      read_ack => Block4_starting_pipe_read_ack,
      read_data => Block4_starting_pipe_read_data,
      write_req => Block4_starting_pipe_write_req,
      write_ack => Block4_starting_pipe_write_ack,
      write_data => Block4_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block5_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block5_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block5_complete_pipe_read_req,
      read_ack => Block5_complete_pipe_read_ack,
      read_data => Block5_complete_pipe_read_data,
      write_req => Block5_complete_pipe_write_req,
      write_ack => Block5_complete_pipe_write_ack,
      write_data => Block5_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block5_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block5_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block5_starting_pipe_read_req,
      read_ack => Block5_starting_pipe_read_ack,
      read_data => Block5_starting_pipe_read_data,
      write_req => Block5_starting_pipe_write_req,
      write_ack => Block5_starting_pipe_write_ack,
      write_data => Block5_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block6_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block6_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block6_complete_pipe_read_req,
      read_ack => Block6_complete_pipe_read_ack,
      read_data => Block6_complete_pipe_read_data,
      write_req => Block6_complete_pipe_write_req,
      write_ack => Block6_complete_pipe_write_ack,
      write_data => Block6_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block6_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block6_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block6_starting_pipe_read_req,
      read_ack => Block6_starting_pipe_read_ack,
      read_data => Block6_starting_pipe_read_data,
      write_req => Block6_starting_pipe_write_req,
      write_ack => Block6_starting_pipe_write_ack,
      write_data => Block6_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block7_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block7_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block7_complete_pipe_read_req,
      read_ack => Block7_complete_pipe_read_ack,
      read_data => Block7_complete_pipe_read_data,
      write_req => Block7_complete_pipe_write_req,
      write_ack => Block7_complete_pipe_write_ack,
      write_data => Block7_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block7_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block7_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block7_starting_pipe_read_req,
      read_ack => Block7_starting_pipe_read_ack,
      read_data => Block7_starting_pipe_read_data,
      write_req => Block7_starting_pipe_write_req,
      write_ack => Block7_starting_pipe_write_ack,
      write_data => Block7_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 8,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 19,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 8,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 19,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyROM_memory_space_2: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
